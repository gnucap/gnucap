
.subckt grids top1 top100 bot50
.parameter r=1
.parameter l=1e-6
.parameter c=1e-9
Rtop_1_2 top1 top2 {r}
Ltop_1_2 top1 top2 {l}
Rbot_1_2 bot1 bot2 {r}
Lbot_1_2 bot1 bot2 {l}
Rtop_1_11 top1 top11 {r}
Ltop_1_11 top1 top11 {l}
Rbot_1_11 bot1 bot11 {r}
Lbot_1_11 bot1 bot11 {l}
C1 top1 bot1 {c}
Rtop_2_3 top2 top3 {r}
Ltop_2_3 top2 top3 {l}
Rbot_2_3 bot2 bot3 {r}
Lbot_2_3 bot2 bot3 {l}
Rtop_2_12 top2 top12 {r}
Ltop_2_12 top2 top12 {l}
Rbot_2_12 bot2 bot12 {r}
Lbot_2_12 bot2 bot12 {l}
C2 top2 bot2 {c}
Rtop_3_4 top3 top4 {r}
Ltop_3_4 top3 top4 {l}
Rbot_3_4 bot3 bot4 {r}
Lbot_3_4 bot3 bot4 {l}
Rtop_3_13 top3 top13 {r}
Ltop_3_13 top3 top13 {l}
Rbot_3_13 bot3 bot13 {r}
Lbot_3_13 bot3 bot13 {l}
C3 top3 bot3 {c}
Rtop_4_5 top4 top5 {r}
Ltop_4_5 top4 top5 {l}
Rbot_4_5 bot4 bot5 {r}
Lbot_4_5 bot4 bot5 {l}
Rtop_4_14 top4 top14 {r}
Ltop_4_14 top4 top14 {l}
Rbot_4_14 bot4 bot14 {r}
Lbot_4_14 bot4 bot14 {l}
C4 top4 bot4 {c}
Rtop_5_6 top5 top6 {r}
Ltop_5_6 top5 top6 {l}
Rbot_5_6 bot5 bot6 {r}
Lbot_5_6 bot5 bot6 {l}
Rtop_5_15 top5 top15 {r}
Ltop_5_15 top5 top15 {l}
Rbot_5_15 bot5 bot15 {r}
Lbot_5_15 bot5 bot15 {l}
C5 top5 bot5 {c}
Rtop_6_7 top6 top7 {r}
Ltop_6_7 top6 top7 {l}
Rbot_6_7 bot6 bot7 {r}
Lbot_6_7 bot6 bot7 {l}
Rtop_6_16 top6 top16 {r}
Ltop_6_16 top6 top16 {l}
Rbot_6_16 bot6 bot16 {r}
Lbot_6_16 bot6 bot16 {l}
C6 top6 bot6 {c}
Rtop_7_8 top7 top8 {r}
Ltop_7_8 top7 top8 {l}
Rbot_7_8 bot7 bot8 {r}
Lbot_7_8 bot7 bot8 {l}
Rtop_7_17 top7 top17 {r}
Ltop_7_17 top7 top17 {l}
Rbot_7_17 bot7 bot17 {r}
Lbot_7_17 bot7 bot17 {l}
C7 top7 bot7 {c}
Rtop_8_9 top8 top9 {r}
Ltop_8_9 top8 top9 {l}
Rbot_8_9 bot8 bot9 {r}
Lbot_8_9 bot8 bot9 {l}
Rtop_8_18 top8 top18 {r}
Ltop_8_18 top8 top18 {l}
Rbot_8_18 bot8 bot18 {r}
Lbot_8_18 bot8 bot18 {l}
C8 top8 bot8 {c}
Rtop_9_10 top9 top10 {r}
Ltop_9_10 top9 top10 {l}
Rbot_9_10 bot9 bot10 {r}
Lbot_9_10 bot9 bot10 {l}
Rtop_9_19 top9 top19 {r}
Ltop_9_19 top9 top19 {l}
Rbot_9_19 bot9 bot19 {r}
Lbot_9_19 bot9 bot19 {l}
C9 top9 bot9 {c}
Rtop_10_20 top10 top20 {r}
Ltop_10_20 top10 top20 {l}
Rbot_10_20 bot10 bot20 {r}
Lbot_10_20 bot10 bot20 {l}
C10 top10 bot10 {c}
Rtop_11_12 top11 top12 {r}
Ltop_11_12 top11 top12 {l}
Rbot_11_12 bot11 bot12 {r}
Lbot_11_12 bot11 bot12 {l}
Rtop_11_21 top11 top21 {r}
Ltop_11_21 top11 top21 {l}
Rbot_11_21 bot11 bot21 {r}
Lbot_11_21 bot11 bot21 {l}
C11 top11 bot11 {c}
Rtop_12_13 top12 top13 {r}
Ltop_12_13 top12 top13 {l}
Rbot_12_13 bot12 bot13 {r}
Lbot_12_13 bot12 bot13 {l}
Rtop_12_22 top12 top22 {r}
Ltop_12_22 top12 top22 {l}
Rbot_12_22 bot12 bot22 {r}
Lbot_12_22 bot12 bot22 {l}
C12 top12 bot12 {c}
Rtop_13_14 top13 top14 {r}
Ltop_13_14 top13 top14 {l}
Rbot_13_14 bot13 bot14 {r}
Lbot_13_14 bot13 bot14 {l}
Rtop_13_23 top13 top23 {r}
Ltop_13_23 top13 top23 {l}
Rbot_13_23 bot13 bot23 {r}
Lbot_13_23 bot13 bot23 {l}
C13 top13 bot13 {c}
Rtop_14_15 top14 top15 {r}
Ltop_14_15 top14 top15 {l}
Rbot_14_15 bot14 bot15 {r}
Lbot_14_15 bot14 bot15 {l}
Rtop_14_24 top14 top24 {r}
Ltop_14_24 top14 top24 {l}
Rbot_14_24 bot14 bot24 {r}
Lbot_14_24 bot14 bot24 {l}
C14 top14 bot14 {c}
Rtop_15_16 top15 top16 {r}
Ltop_15_16 top15 top16 {l}
Rbot_15_16 bot15 bot16 {r}
Lbot_15_16 bot15 bot16 {l}
Rtop_15_25 top15 top25 {r}
Ltop_15_25 top15 top25 {l}
Rbot_15_25 bot15 bot25 {r}
Lbot_15_25 bot15 bot25 {l}
C15 top15 bot15 {c}
Rtop_16_17 top16 top17 {r}
Ltop_16_17 top16 top17 {l}
Rbot_16_17 bot16 bot17 {r}
Lbot_16_17 bot16 bot17 {l}
Rtop_16_26 top16 top26 {r}
Ltop_16_26 top16 top26 {l}
Rbot_16_26 bot16 bot26 {r}
Lbot_16_26 bot16 bot26 {l}
C16 top16 bot16 {c}
Rtop_17_18 top17 top18 {r}
Ltop_17_18 top17 top18 {l}
Rbot_17_18 bot17 bot18 {r}
Lbot_17_18 bot17 bot18 {l}
Rtop_17_27 top17 top27 {r}
Ltop_17_27 top17 top27 {l}
Rbot_17_27 bot17 bot27 {r}
Lbot_17_27 bot17 bot27 {l}
C17 top17 bot17 {c}
Rtop_18_19 top18 top19 {r}
Ltop_18_19 top18 top19 {l}
Rbot_18_19 bot18 bot19 {r}
Lbot_18_19 bot18 bot19 {l}
Rtop_18_28 top18 top28 {r}
Ltop_18_28 top18 top28 {l}
Rbot_18_28 bot18 bot28 {r}
Lbot_18_28 bot18 bot28 {l}
C18 top18 bot18 {c}
Rtop_19_20 top19 top20 {r}
Ltop_19_20 top19 top20 {l}
Rbot_19_20 bot19 bot20 {r}
Lbot_19_20 bot19 bot20 {l}
Rtop_19_29 top19 top29 {r}
Ltop_19_29 top19 top29 {l}
Rbot_19_29 bot19 bot29 {r}
Lbot_19_29 bot19 bot29 {l}
C19 top19 bot19 {c}
Rtop_20_30 top20 top30 {r}
Ltop_20_30 top20 top30 {l}
Rbot_20_30 bot20 bot30 {r}
Lbot_20_30 bot20 bot30 {l}
C20 top20 bot20 {c}
Rtop_21_22 top21 top22 {r}
Ltop_21_22 top21 top22 {l}
Rbot_21_22 bot21 bot22 {r}
Lbot_21_22 bot21 bot22 {l}
Rtop_21_31 top21 top31 {r}
Ltop_21_31 top21 top31 {l}
Rbot_21_31 bot21 bot31 {r}
Lbot_21_31 bot21 bot31 {l}
C21 top21 bot21 {c}
Rtop_22_23 top22 top23 {r}
Ltop_22_23 top22 top23 {l}
Rbot_22_23 bot22 bot23 {r}
Lbot_22_23 bot22 bot23 {l}
Rtop_22_32 top22 top32 {r}
Ltop_22_32 top22 top32 {l}
Rbot_22_32 bot22 bot32 {r}
Lbot_22_32 bot22 bot32 {l}
C22 top22 bot22 {c}
Rtop_23_24 top23 top24 {r}
Ltop_23_24 top23 top24 {l}
Rbot_23_24 bot23 bot24 {r}
Lbot_23_24 bot23 bot24 {l}
Rtop_23_33 top23 top33 {r}
Ltop_23_33 top23 top33 {l}
Rbot_23_33 bot23 bot33 {r}
Lbot_23_33 bot23 bot33 {l}
C23 top23 bot23 {c}
Rtop_24_25 top24 top25 {r}
Ltop_24_25 top24 top25 {l}
Rbot_24_25 bot24 bot25 {r}
Lbot_24_25 bot24 bot25 {l}
Rtop_24_34 top24 top34 {r}
Ltop_24_34 top24 top34 {l}
Rbot_24_34 bot24 bot34 {r}
Lbot_24_34 bot24 bot34 {l}
C24 top24 bot24 {c}
Rtop_25_26 top25 top26 {r}
Ltop_25_26 top25 top26 {l}
Rbot_25_26 bot25 bot26 {r}
Lbot_25_26 bot25 bot26 {l}
Rtop_25_35 top25 top35 {r}
Ltop_25_35 top25 top35 {l}
Rbot_25_35 bot25 bot35 {r}
Lbot_25_35 bot25 bot35 {l}
C25 top25 bot25 {c}
Rtop_26_27 top26 top27 {r}
Ltop_26_27 top26 top27 {l}
Rbot_26_27 bot26 bot27 {r}
Lbot_26_27 bot26 bot27 {l}
Rtop_26_36 top26 top36 {r}
Ltop_26_36 top26 top36 {l}
Rbot_26_36 bot26 bot36 {r}
Lbot_26_36 bot26 bot36 {l}
C26 top26 bot26 {c}
Rtop_27_28 top27 top28 {r}
Ltop_27_28 top27 top28 {l}
Rbot_27_28 bot27 bot28 {r}
Lbot_27_28 bot27 bot28 {l}
Rtop_27_37 top27 top37 {r}
Ltop_27_37 top27 top37 {l}
Rbot_27_37 bot27 bot37 {r}
Lbot_27_37 bot27 bot37 {l}
C27 top27 bot27 {c}
Rtop_28_29 top28 top29 {r}
Ltop_28_29 top28 top29 {l}
Rbot_28_29 bot28 bot29 {r}
Lbot_28_29 bot28 bot29 {l}
Rtop_28_38 top28 top38 {r}
Ltop_28_38 top28 top38 {l}
Rbot_28_38 bot28 bot38 {r}
Lbot_28_38 bot28 bot38 {l}
C28 top28 bot28 {c}
Rtop_29_30 top29 top30 {r}
Ltop_29_30 top29 top30 {l}
Rbot_29_30 bot29 bot30 {r}
Lbot_29_30 bot29 bot30 {l}
Rtop_29_39 top29 top39 {r}
Ltop_29_39 top29 top39 {l}
Rbot_29_39 bot29 bot39 {r}
Lbot_29_39 bot29 bot39 {l}
C29 top29 bot29 {c}
Rtop_30_40 top30 top40 {r}
Ltop_30_40 top30 top40 {l}
Rbot_30_40 bot30 bot40 {r}
Lbot_30_40 bot30 bot40 {l}
C30 top30 bot30 {c}
Rtop_31_32 top31 top32 {r}
Ltop_31_32 top31 top32 {l}
Rbot_31_32 bot31 bot32 {r}
Lbot_31_32 bot31 bot32 {l}
Rtop_31_41 top31 top41 {r}
Ltop_31_41 top31 top41 {l}
Rbot_31_41 bot31 bot41 {r}
Lbot_31_41 bot31 bot41 {l}
C31 top31 bot31 {c}
Rtop_32_33 top32 top33 {r}
Ltop_32_33 top32 top33 {l}
Rbot_32_33 bot32 bot33 {r}
Lbot_32_33 bot32 bot33 {l}
Rtop_32_42 top32 top42 {r}
Ltop_32_42 top32 top42 {l}
Rbot_32_42 bot32 bot42 {r}
Lbot_32_42 bot32 bot42 {l}
C32 top32 bot32 {c}
Rtop_33_34 top33 top34 {r}
Ltop_33_34 top33 top34 {l}
Rbot_33_34 bot33 bot34 {r}
Lbot_33_34 bot33 bot34 {l}
Rtop_33_43 top33 top43 {r}
Ltop_33_43 top33 top43 {l}
Rbot_33_43 bot33 bot43 {r}
Lbot_33_43 bot33 bot43 {l}
C33 top33 bot33 {c}
Rtop_34_35 top34 top35 {r}
Ltop_34_35 top34 top35 {l}
Rbot_34_35 bot34 bot35 {r}
Lbot_34_35 bot34 bot35 {l}
Rtop_34_44 top34 top44 {r}
Ltop_34_44 top34 top44 {l}
Rbot_34_44 bot34 bot44 {r}
Lbot_34_44 bot34 bot44 {l}
C34 top34 bot34 {c}
Rtop_35_36 top35 top36 {r}
Ltop_35_36 top35 top36 {l}
Rbot_35_36 bot35 bot36 {r}
Lbot_35_36 bot35 bot36 {l}
Rtop_35_45 top35 top45 {r}
Ltop_35_45 top35 top45 {l}
Rbot_35_45 bot35 bot45 {r}
Lbot_35_45 bot35 bot45 {l}
C35 top35 bot35 {c}
Rtop_36_37 top36 top37 {r}
Ltop_36_37 top36 top37 {l}
Rbot_36_37 bot36 bot37 {r}
Lbot_36_37 bot36 bot37 {l}
Rtop_36_46 top36 top46 {r}
Ltop_36_46 top36 top46 {l}
Rbot_36_46 bot36 bot46 {r}
Lbot_36_46 bot36 bot46 {l}
C36 top36 bot36 {c}
Rtop_37_38 top37 top38 {r}
Ltop_37_38 top37 top38 {l}
Rbot_37_38 bot37 bot38 {r}
Lbot_37_38 bot37 bot38 {l}
Rtop_37_47 top37 top47 {r}
Ltop_37_47 top37 top47 {l}
Rbot_37_47 bot37 bot47 {r}
Lbot_37_47 bot37 bot47 {l}
C37 top37 bot37 {c}
Rtop_38_39 top38 top39 {r}
Ltop_38_39 top38 top39 {l}
Rbot_38_39 bot38 bot39 {r}
Lbot_38_39 bot38 bot39 {l}
Rtop_38_48 top38 top48 {r}
Ltop_38_48 top38 top48 {l}
Rbot_38_48 bot38 bot48 {r}
Lbot_38_48 bot38 bot48 {l}
C38 top38 bot38 {c}
Rtop_39_40 top39 top40 {r}
Ltop_39_40 top39 top40 {l}
Rbot_39_40 bot39 bot40 {r}
Lbot_39_40 bot39 bot40 {l}
Rtop_39_49 top39 top49 {r}
Ltop_39_49 top39 top49 {l}
Rbot_39_49 bot39 bot49 {r}
Lbot_39_49 bot39 bot49 {l}
C39 top39 bot39 {c}
Rtop_40_50 top40 top50 {r}
Ltop_40_50 top40 top50 {l}
Rbot_40_50 bot40 bot50 {r}
Lbot_40_50 bot40 bot50 {l}
C40 top40 bot40 {c}
Rtop_41_42 top41 top42 {r}
Ltop_41_42 top41 top42 {l}
Rbot_41_42 bot41 bot42 {r}
Lbot_41_42 bot41 bot42 {l}
Rtop_41_51 top41 top51 {r}
Ltop_41_51 top41 top51 {l}
Rbot_41_51 bot41 bot51 {r}
Lbot_41_51 bot41 bot51 {l}
C41 top41 bot41 {c}
Rtop_42_43 top42 top43 {r}
Ltop_42_43 top42 top43 {l}
Rbot_42_43 bot42 bot43 {r}
Lbot_42_43 bot42 bot43 {l}
Rtop_42_52 top42 top52 {r}
Ltop_42_52 top42 top52 {l}
Rbot_42_52 bot42 bot52 {r}
Lbot_42_52 bot42 bot52 {l}
C42 top42 bot42 {c}
Rtop_43_44 top43 top44 {r}
Ltop_43_44 top43 top44 {l}
Rbot_43_44 bot43 bot44 {r}
Lbot_43_44 bot43 bot44 {l}
Rtop_43_53 top43 top53 {r}
Ltop_43_53 top43 top53 {l}
Rbot_43_53 bot43 bot53 {r}
Lbot_43_53 bot43 bot53 {l}
C43 top43 bot43 {c}
Rtop_44_45 top44 top45 {r}
Ltop_44_45 top44 top45 {l}
Rbot_44_45 bot44 bot45 {r}
Lbot_44_45 bot44 bot45 {l}
Rtop_44_54 top44 top54 {r}
Ltop_44_54 top44 top54 {l}
Rbot_44_54 bot44 bot54 {r}
Lbot_44_54 bot44 bot54 {l}
C44 top44 bot44 {c}
Rtop_45_46 top45 top46 {r}
Ltop_45_46 top45 top46 {l}
Rbot_45_46 bot45 bot46 {r}
Lbot_45_46 bot45 bot46 {l}
Rtop_45_55 top45 top55 {r}
Ltop_45_55 top45 top55 {l}
Rbot_45_55 bot45 bot55 {r}
Lbot_45_55 bot45 bot55 {l}
C45 top45 bot45 {c}
Rtop_46_47 top46 top47 {r}
Ltop_46_47 top46 top47 {l}
Rbot_46_47 bot46 bot47 {r}
Lbot_46_47 bot46 bot47 {l}
Rtop_46_56 top46 top56 {r}
Ltop_46_56 top46 top56 {l}
Rbot_46_56 bot46 bot56 {r}
Lbot_46_56 bot46 bot56 {l}
C46 top46 bot46 {c}
Rtop_47_48 top47 top48 {r}
Ltop_47_48 top47 top48 {l}
Rbot_47_48 bot47 bot48 {r}
Lbot_47_48 bot47 bot48 {l}
Rtop_47_57 top47 top57 {r}
Ltop_47_57 top47 top57 {l}
Rbot_47_57 bot47 bot57 {r}
Lbot_47_57 bot47 bot57 {l}
C47 top47 bot47 {c}
Rtop_48_49 top48 top49 {r}
Ltop_48_49 top48 top49 {l}
Rbot_48_49 bot48 bot49 {r}
Lbot_48_49 bot48 bot49 {l}
Rtop_48_58 top48 top58 {r}
Ltop_48_58 top48 top58 {l}
Rbot_48_58 bot48 bot58 {r}
Lbot_48_58 bot48 bot58 {l}
C48 top48 bot48 {c}
Rtop_49_50 top49 top50 {r}
Ltop_49_50 top49 top50 {l}
Rbot_49_50 bot49 bot50 {r}
Lbot_49_50 bot49 bot50 {l}
Rtop_49_59 top49 top59 {r}
Ltop_49_59 top49 top59 {l}
Rbot_49_59 bot49 bot59 {r}
Lbot_49_59 bot49 bot59 {l}
C49 top49 bot49 {c}
Rtop_50_60 top50 top60 {r}
Ltop_50_60 top50 top60 {l}
Rbot_50_60 bot50 bot60 {r}
Lbot_50_60 bot50 bot60 {l}
C50 top50 bot50 {c}
Rtop_51_52 top51 top52 {r}
Ltop_51_52 top51 top52 {l}
Rbot_51_52 bot51 bot52 {r}
Lbot_51_52 bot51 bot52 {l}
Rtop_51_61 top51 top61 {r}
Ltop_51_61 top51 top61 {l}
Rbot_51_61 bot51 bot61 {r}
Lbot_51_61 bot51 bot61 {l}
C51 top51 bot51 {c}
Rtop_52_53 top52 top53 {r}
Ltop_52_53 top52 top53 {l}
Rbot_52_53 bot52 bot53 {r}
Lbot_52_53 bot52 bot53 {l}
Rtop_52_62 top52 top62 {r}
Ltop_52_62 top52 top62 {l}
Rbot_52_62 bot52 bot62 {r}
Lbot_52_62 bot52 bot62 {l}
C52 top52 bot52 {c}
Rtop_53_54 top53 top54 {r}
Ltop_53_54 top53 top54 {l}
Rbot_53_54 bot53 bot54 {r}
Lbot_53_54 bot53 bot54 {l}
Rtop_53_63 top53 top63 {r}
Ltop_53_63 top53 top63 {l}
Rbot_53_63 bot53 bot63 {r}
Lbot_53_63 bot53 bot63 {l}
C53 top53 bot53 {c}
Rtop_54_55 top54 top55 {r}
Ltop_54_55 top54 top55 {l}
Rbot_54_55 bot54 bot55 {r}
Lbot_54_55 bot54 bot55 {l}
Rtop_54_64 top54 top64 {r}
Ltop_54_64 top54 top64 {l}
Rbot_54_64 bot54 bot64 {r}
Lbot_54_64 bot54 bot64 {l}
C54 top54 bot54 {c}
Rtop_55_56 top55 top56 {r}
Ltop_55_56 top55 top56 {l}
Rbot_55_56 bot55 bot56 {r}
Lbot_55_56 bot55 bot56 {l}
Rtop_55_65 top55 top65 {r}
Ltop_55_65 top55 top65 {l}
Rbot_55_65 bot55 bot65 {r}
Lbot_55_65 bot55 bot65 {l}
C55 top55 bot55 {c}
Rtop_56_57 top56 top57 {r}
Ltop_56_57 top56 top57 {l}
Rbot_56_57 bot56 bot57 {r}
Lbot_56_57 bot56 bot57 {l}
Rtop_56_66 top56 top66 {r}
Ltop_56_66 top56 top66 {l}
Rbot_56_66 bot56 bot66 {r}
Lbot_56_66 bot56 bot66 {l}
C56 top56 bot56 {c}
Rtop_57_58 top57 top58 {r}
Ltop_57_58 top57 top58 {l}
Rbot_57_58 bot57 bot58 {r}
Lbot_57_58 bot57 bot58 {l}
Rtop_57_67 top57 top67 {r}
Ltop_57_67 top57 top67 {l}
Rbot_57_67 bot57 bot67 {r}
Lbot_57_67 bot57 bot67 {l}
C57 top57 bot57 {c}
Rtop_58_59 top58 top59 {r}
Ltop_58_59 top58 top59 {l}
Rbot_58_59 bot58 bot59 {r}
Lbot_58_59 bot58 bot59 {l}
Rtop_58_68 top58 top68 {r}
Ltop_58_68 top58 top68 {l}
Rbot_58_68 bot58 bot68 {r}
Lbot_58_68 bot58 bot68 {l}
C58 top58 bot58 {c}
Rtop_59_60 top59 top60 {r}
Ltop_59_60 top59 top60 {l}
Rbot_59_60 bot59 bot60 {r}
Lbot_59_60 bot59 bot60 {l}
Rtop_59_69 top59 top69 {r}
Ltop_59_69 top59 top69 {l}
Rbot_59_69 bot59 bot69 {r}
Lbot_59_69 bot59 bot69 {l}
C59 top59 bot59 {c}
Rtop_60_70 top60 top70 {r}
Ltop_60_70 top60 top70 {l}
Rbot_60_70 bot60 bot70 {r}
Lbot_60_70 bot60 bot70 {l}
C60 top60 bot60 {c}
Rtop_61_62 top61 top62 {r}
Ltop_61_62 top61 top62 {l}
Rbot_61_62 bot61 bot62 {r}
Lbot_61_62 bot61 bot62 {l}
Rtop_61_71 top61 top71 {r}
Ltop_61_71 top61 top71 {l}
Rbot_61_71 bot61 bot71 {r}
Lbot_61_71 bot61 bot71 {l}
C61 top61 bot61 {c}
Rtop_62_63 top62 top63 {r}
Ltop_62_63 top62 top63 {l}
Rbot_62_63 bot62 bot63 {r}
Lbot_62_63 bot62 bot63 {l}
Rtop_62_72 top62 top72 {r}
Ltop_62_72 top62 top72 {l}
Rbot_62_72 bot62 bot72 {r}
Lbot_62_72 bot62 bot72 {l}
C62 top62 bot62 {c}
Rtop_63_64 top63 top64 {r}
Ltop_63_64 top63 top64 {l}
Rbot_63_64 bot63 bot64 {r}
Lbot_63_64 bot63 bot64 {l}
Rtop_63_73 top63 top73 {r}
Ltop_63_73 top63 top73 {l}
Rbot_63_73 bot63 bot73 {r}
Lbot_63_73 bot63 bot73 {l}
C63 top63 bot63 {c}
Rtop_64_65 top64 top65 {r}
Ltop_64_65 top64 top65 {l}
Rbot_64_65 bot64 bot65 {r}
Lbot_64_65 bot64 bot65 {l}
Rtop_64_74 top64 top74 {r}
Ltop_64_74 top64 top74 {l}
Rbot_64_74 bot64 bot74 {r}
Lbot_64_74 bot64 bot74 {l}
C64 top64 bot64 {c}
Rtop_65_66 top65 top66 {r}
Ltop_65_66 top65 top66 {l}
Rbot_65_66 bot65 bot66 {r}
Lbot_65_66 bot65 bot66 {l}
Rtop_65_75 top65 top75 {r}
Ltop_65_75 top65 top75 {l}
Rbot_65_75 bot65 bot75 {r}
Lbot_65_75 bot65 bot75 {l}
C65 top65 bot65 {c}
Rtop_66_67 top66 top67 {r}
Ltop_66_67 top66 top67 {l}
Rbot_66_67 bot66 bot67 {r}
Lbot_66_67 bot66 bot67 {l}
Rtop_66_76 top66 top76 {r}
Ltop_66_76 top66 top76 {l}
Rbot_66_76 bot66 bot76 {r}
Lbot_66_76 bot66 bot76 {l}
C66 top66 bot66 {c}
Rtop_67_68 top67 top68 {r}
Ltop_67_68 top67 top68 {l}
Rbot_67_68 bot67 bot68 {r}
Lbot_67_68 bot67 bot68 {l}
Rtop_67_77 top67 top77 {r}
Ltop_67_77 top67 top77 {l}
Rbot_67_77 bot67 bot77 {r}
Lbot_67_77 bot67 bot77 {l}
C67 top67 bot67 {c}
Rtop_68_69 top68 top69 {r}
Ltop_68_69 top68 top69 {l}
Rbot_68_69 bot68 bot69 {r}
Lbot_68_69 bot68 bot69 {l}
Rtop_68_78 top68 top78 {r}
Ltop_68_78 top68 top78 {l}
Rbot_68_78 bot68 bot78 {r}
Lbot_68_78 bot68 bot78 {l}
C68 top68 bot68 {c}
Rtop_69_70 top69 top70 {r}
Ltop_69_70 top69 top70 {l}
Rbot_69_70 bot69 bot70 {r}
Lbot_69_70 bot69 bot70 {l}
Rtop_69_79 top69 top79 {r}
Ltop_69_79 top69 top79 {l}
Rbot_69_79 bot69 bot79 {r}
Lbot_69_79 bot69 bot79 {l}
C69 top69 bot69 {c}
Rtop_70_80 top70 top80 {r}
Ltop_70_80 top70 top80 {l}
Rbot_70_80 bot70 bot80 {r}
Lbot_70_80 bot70 bot80 {l}
C70 top70 bot70 {c}
Rtop_71_72 top71 top72 {r}
Ltop_71_72 top71 top72 {l}
Rbot_71_72 bot71 bot72 {r}
Lbot_71_72 bot71 bot72 {l}
Rtop_71_81 top71 top81 {r}
Ltop_71_81 top71 top81 {l}
Rbot_71_81 bot71 bot81 {r}
Lbot_71_81 bot71 bot81 {l}
C71 top71 bot71 {c}
Rtop_72_73 top72 top73 {r}
Ltop_72_73 top72 top73 {l}
Rbot_72_73 bot72 bot73 {r}
Lbot_72_73 bot72 bot73 {l}
Rtop_72_82 top72 top82 {r}
Ltop_72_82 top72 top82 {l}
Rbot_72_82 bot72 bot82 {r}
Lbot_72_82 bot72 bot82 {l}
C72 top72 bot72 {c}
Rtop_73_74 top73 top74 {r}
Ltop_73_74 top73 top74 {l}
Rbot_73_74 bot73 bot74 {r}
Lbot_73_74 bot73 bot74 {l}
Rtop_73_83 top73 top83 {r}
Ltop_73_83 top73 top83 {l}
Rbot_73_83 bot73 bot83 {r}
Lbot_73_83 bot73 bot83 {l}
C73 top73 bot73 {c}
Rtop_74_75 top74 top75 {r}
Ltop_74_75 top74 top75 {l}
Rbot_74_75 bot74 bot75 {r}
Lbot_74_75 bot74 bot75 {l}
Rtop_74_84 top74 top84 {r}
Ltop_74_84 top74 top84 {l}
Rbot_74_84 bot74 bot84 {r}
Lbot_74_84 bot74 bot84 {l}
C74 top74 bot74 {c}
Rtop_75_76 top75 top76 {r}
Ltop_75_76 top75 top76 {l}
Rbot_75_76 bot75 bot76 {r}
Lbot_75_76 bot75 bot76 {l}
Rtop_75_85 top75 top85 {r}
Ltop_75_85 top75 top85 {l}
Rbot_75_85 bot75 bot85 {r}
Lbot_75_85 bot75 bot85 {l}
C75 top75 bot75 {c}
Rtop_76_77 top76 top77 {r}
Ltop_76_77 top76 top77 {l}
Rbot_76_77 bot76 bot77 {r}
Lbot_76_77 bot76 bot77 {l}
Rtop_76_86 top76 top86 {r}
Ltop_76_86 top76 top86 {l}
Rbot_76_86 bot76 bot86 {r}
Lbot_76_86 bot76 bot86 {l}
C76 top76 bot76 {c}
Rtop_77_78 top77 top78 {r}
Ltop_77_78 top77 top78 {l}
Rbot_77_78 bot77 bot78 {r}
Lbot_77_78 bot77 bot78 {l}
Rtop_77_87 top77 top87 {r}
Ltop_77_87 top77 top87 {l}
Rbot_77_87 bot77 bot87 {r}
Lbot_77_87 bot77 bot87 {l}
C77 top77 bot77 {c}
Rtop_78_79 top78 top79 {r}
Ltop_78_79 top78 top79 {l}
Rbot_78_79 bot78 bot79 {r}
Lbot_78_79 bot78 bot79 {l}
Rtop_78_88 top78 top88 {r}
Ltop_78_88 top78 top88 {l}
Rbot_78_88 bot78 bot88 {r}
Lbot_78_88 bot78 bot88 {l}
C78 top78 bot78 {c}
Rtop_79_80 top79 top80 {r}
Ltop_79_80 top79 top80 {l}
Rbot_79_80 bot79 bot80 {r}
Lbot_79_80 bot79 bot80 {l}
Rtop_79_89 top79 top89 {r}
Ltop_79_89 top79 top89 {l}
Rbot_79_89 bot79 bot89 {r}
Lbot_79_89 bot79 bot89 {l}
C79 top79 bot79 {c}
Rtop_80_90 top80 top90 {r}
Ltop_80_90 top80 top90 {l}
Rbot_80_90 bot80 bot90 {r}
Lbot_80_90 bot80 bot90 {l}
C80 top80 bot80 {c}
Rtop_81_82 top81 top82 {r}
Ltop_81_82 top81 top82 {l}
Rbot_81_82 bot81 bot82 {r}
Lbot_81_82 bot81 bot82 {l}
Rtop_81_91 top81 top91 {r}
Ltop_81_91 top81 top91 {l}
Rbot_81_91 bot81 bot91 {r}
Lbot_81_91 bot81 bot91 {l}
C81 top81 bot81 {c}
Rtop_82_83 top82 top83 {r}
Ltop_82_83 top82 top83 {l}
Rbot_82_83 bot82 bot83 {r}
Lbot_82_83 bot82 bot83 {l}
Rtop_82_92 top82 top92 {r}
Ltop_82_92 top82 top92 {l}
Rbot_82_92 bot82 bot92 {r}
Lbot_82_92 bot82 bot92 {l}
C82 top82 bot82 {c}
Rtop_83_84 top83 top84 {r}
Ltop_83_84 top83 top84 {l}
Rbot_83_84 bot83 bot84 {r}
Lbot_83_84 bot83 bot84 {l}
Rtop_83_93 top83 top93 {r}
Ltop_83_93 top83 top93 {l}
Rbot_83_93 bot83 bot93 {r}
Lbot_83_93 bot83 bot93 {l}
C83 top83 bot83 {c}
Rtop_84_85 top84 top85 {r}
Ltop_84_85 top84 top85 {l}
Rbot_84_85 bot84 bot85 {r}
Lbot_84_85 bot84 bot85 {l}
Rtop_84_94 top84 top94 {r}
Ltop_84_94 top84 top94 {l}
Rbot_84_94 bot84 bot94 {r}
Lbot_84_94 bot84 bot94 {l}
C84 top84 bot84 {c}
Rtop_85_86 top85 top86 {r}
Ltop_85_86 top85 top86 {l}
Rbot_85_86 bot85 bot86 {r}
Lbot_85_86 bot85 bot86 {l}
Rtop_85_95 top85 top95 {r}
Ltop_85_95 top85 top95 {l}
Rbot_85_95 bot85 bot95 {r}
Lbot_85_95 bot85 bot95 {l}
C85 top85 bot85 {c}
Rtop_86_87 top86 top87 {r}
Ltop_86_87 top86 top87 {l}
Rbot_86_87 bot86 bot87 {r}
Lbot_86_87 bot86 bot87 {l}
Rtop_86_96 top86 top96 {r}
Ltop_86_96 top86 top96 {l}
Rbot_86_96 bot86 bot96 {r}
Lbot_86_96 bot86 bot96 {l}
C86 top86 bot86 {c}
Rtop_87_88 top87 top88 {r}
Ltop_87_88 top87 top88 {l}
Rbot_87_88 bot87 bot88 {r}
Lbot_87_88 bot87 bot88 {l}
Rtop_87_97 top87 top97 {r}
Ltop_87_97 top87 top97 {l}
Rbot_87_97 bot87 bot97 {r}
Lbot_87_97 bot87 bot97 {l}
C87 top87 bot87 {c}
Rtop_88_89 top88 top89 {r}
Ltop_88_89 top88 top89 {l}
Rbot_88_89 bot88 bot89 {r}
Lbot_88_89 bot88 bot89 {l}
Rtop_88_98 top88 top98 {r}
Ltop_88_98 top88 top98 {l}
Rbot_88_98 bot88 bot98 {r}
Lbot_88_98 bot88 bot98 {l}
C88 top88 bot88 {c}
Rtop_89_90 top89 top90 {r}
Ltop_89_90 top89 top90 {l}
Rbot_89_90 bot89 bot90 {r}
Lbot_89_90 bot89 bot90 {l}
Rtop_89_99 top89 top99 {r}
Ltop_89_99 top89 top99 {l}
Rbot_89_99 bot89 bot99 {r}
Lbot_89_99 bot89 bot99 {l}
C89 top89 bot89 {c}
Rtop_90_100 top90 top100 {r}
Ltop_90_100 top90 top100 {l}
Rbot_90_100 bot90 bot100 {r}
Lbot_90_100 bot90 bot100 {l}
C90 top90 bot90 {c}
Rtop_91_92 top91 top92 {r}
Ltop_91_92 top91 top92 {l}
Rbot_91_92 bot91 bot92 {r}
Lbot_91_92 bot91 bot92 {l}
C91 top91 bot91 {c}
Rtop_92_93 top92 top93 {r}
Ltop_92_93 top92 top93 {l}
Rbot_92_93 bot92 bot93 {r}
Lbot_92_93 bot92 bot93 {l}
C92 top92 bot92 {c}
Rtop_93_94 top93 top94 {r}
Ltop_93_94 top93 top94 {l}
Rbot_93_94 bot93 bot94 {r}
Lbot_93_94 bot93 bot94 {l}
C93 top93 bot93 {c}
Rtop_94_95 top94 top95 {r}
Ltop_94_95 top94 top95 {l}
Rbot_94_95 bot94 bot95 {r}
Lbot_94_95 bot94 bot95 {l}
C94 top94 bot94 {c}
Rtop_95_96 top95 top96 {r}
Ltop_95_96 top95 top96 {l}
Rbot_95_96 bot95 bot96 {r}
Lbot_95_96 bot95 bot96 {l}
C95 top95 bot95 {c}
Rtop_96_97 top96 top97 {r}
Ltop_96_97 top96 top97 {l}
Rbot_96_97 bot96 bot97 {r}
Lbot_96_97 bot96 bot97 {l}
C96 top96 bot96 {c}
Rtop_97_98 top97 top98 {r}
Ltop_97_98 top97 top98 {l}
Rbot_97_98 bot97 bot98 {r}
Lbot_97_98 bot97 bot98 {l}
C97 top97 bot97 {c}
Rtop_98_99 top98 top99 {r}
Ltop_98_99 top98 top99 {l}
Rbot_98_99 bot98 bot99 {r}
Lbot_98_99 bot98 bot99 {l}
C98 top98 bot98 {c}
Rtop_99_100 top99 top100 {r}
Ltop_99_100 top99 top100 {l}
Rbot_99_100 bot99 bot100 {r}
Lbot_99_100 bot99 bot100 {l}
C99 top99 bot99 {c}
C100 top100 bot100 {c}
.ends

X1 in out 0 grids
v1 in 0 ac 1 dc 0

*>.print ac vr(out) vi(out) vm(out) vp(out)
*>.print op v(out)
*>.op
*>.ac oct 1 1 250k basic

*>.end

* try this with ngspice -b ..
.control
ac oct 1 1 500k
set units = degrees
.endc
.print ac vm(out) vp(out)
