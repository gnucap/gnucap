# expression error
.eval foo(3)
