# expression test
.option list
.param a=9
.eval a
.param b=-8
.eval b
.param c={3*8}
.eval c
.param d={3+8}
.eval d
.param e={3-8}
.eval e
.param f={3/8}
.eval f
.param a1={3==8}
.eval a1
.param b1={3!=8}
.eval b1
.param c1={3<8}
.eval c1
.param d1={3>8}
.eval d1
.param e1={3<=8}
.eval e1
.param f1={3>=8}
.eval f1
.param g1={3||8}
.eval g1
.param h1={3&&8}
.eval h1
.param a2={3==3}
.eval a2
.param b2={3!=3}
.eval b2
.param c2={3<3}
.eval c2
.param d2={3>3}
.eval d2
.param e2={3<=3}
.eval e2
.param f2={3>=3}
.eval f2
.param g2={3||3}
.eval g2
.param h2={3&&3}
.eval h2
.param j1={0||0}
.eval j1
.param j2={0||1}
.eval j2
.param j3={1||0}
.eval j3
.param j4={1||1}
.eval j4
.param k1={0&&0}
.eval k1
.param k2={0&&1}
.eval k2
.param k3={1&&0}
.eval k3
.param k4={1&&1}
.eval k4
