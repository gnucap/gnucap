nmos n gate, saturated
M1   2  2  0  0  cmosn  l= 9.u  w= 9.u  nrd= 1.  nrs= 1. 
Vds   3  0  5.
Rds   2  3  10
.model cmosn  nmos (level=6 tox=1e-7)
.op
.print dc v(1) v(2) v(3) i(vds)
.dc vgs -10 10 1
.end
