' cap with initial condition
c1 1 0 1 ic=3
r1 1 0 1
.list
.print tran v(1)
.tran 1 10 0 uic
.status notime
.end
