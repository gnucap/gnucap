'
V1   2  0  1.
X1   2  1  3 zzz
X2   2  4  5 zzz
.macro zzz  1 2 4
R1   1  2  1.
R2   2  0  1.
R3   2  3  1.
R4   3  0  1.
r5 3 4 1
r6 4 0 1
.eom zzz
.width out=160
.print op v(nodes)
.op
.print op + v(r1.x1) v(r?.x1) v(r2.x?)
.op
.print
.list
.end
