' dc sweep test
v1 1 0 1
v2 2 0 dc 1
v3 3 0 ac 1
r1 1 0 100k
r2 2 0 100k
r3 3 0 100k
.print dc v(1) v(2) v(3)
.dc v1 -2 2 1
.dc v2 -2 2 1
.dc v3 -2 2 1
.end
