'dctran test
V1   1  0  dc generator(1) ac 1
L3   1  2  dc 1. ac 1.
R4   2  0  dc 1. ac 1.
R5   1  3  dc 1. ac 1.
C6   3  0  dc 1. ac 1.
.options short=1p
.print tran iter(0)  v(nodes)
.tran 0 1 .1
.print ac v(nodes)
.ac .001 10 decade
.list
.end
