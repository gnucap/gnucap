# cccs test ref to device that does not exist
i1 1 0 11 ac 11
ri1 1 0 10
e1 2 0 1 0 8
re1 2 0 10
* sense the voltage source (0 volts)
f2 5 0 v3 8
rf2 5 0 10
i2 3 0 11 ac 11
ri2 4 0 10
v2 3 4 0
* sense a live voltage source
f7 7 0 v7 8
rf7 7 0 10
v7 6 0 11 ac 11
rv7 6 0 10
.width out=132
.print op v(1) v(2) v(3) v(4) v(5) v(6) v(7) f(f2) f(f7)
.op
.print tran v(1) v(2) v(3) v(4) v(5) v(6) v(7) f(f2) f(f7)
.tran .05 .1 0
.print ac v(1) v(2) v(3) v(4) v(5) v(6) v(7) f(f2) f(f7)
.ac oct 1 1k 2k
.end
