nonlinear res test

V1 1 0  1.
R1 1 0 PWL 0.1,0 1,1 10,2 100,3
+          1000,4 10000,5 100000,6 1000000,7
+          10000000,8 100000000,9 1000000000,10

.options nopicky
.print dc i(R1) vin(r1) i(v1) iter(0) f(R1) df(R1) in(R1) iof(R1)
.dc v1 0 10 1 loop trace n basic
.stat notime
