100 cascaded NMOS inverters
vd1 2 0 5
md1  3 1 0 0  modeld w=10u l=2u
ml1  2 2 3 0  modell w=2u l=2u
vd2 4 0 5
md2  5 3 0 0  modeld w=10u l=2u
ml2  4 4 5 0  modell w=2u l=2u
vd3 6 0 5
md3  7 5 0 0  modeld w=10u l=2u
ml3  6 6 7 0  modell w=2u l=2u
vd4 8 0 5
md4  9 7 0 0  modeld w=10u l=2u
ml4  8 8 9 0  modell w=2u l=2u
vd5 10 0 5
md5  11 9 0 0  modeld w=10u l=2u
ml5  10 10 11 0  modell w=2u l=2u
vd6 12 0 5
md6  13 11 0 0  modeld w=10u l=2u
ml6  12 12 13 0  modell w=2u l=2u
vd7 14 0 5
md7  15 13 0 0  modeld w=10u l=2u
ml7  14 14 15 0  modell w=2u l=2u
vd8 16 0 5
md8  17 15 0 0  modeld w=10u l=2u
ml8  16 16 17 0  modell w=2u l=2u
vd9 18 0 5
md9  19 17 0 0  modeld w=10u l=2u
ml9  18 18 19 0  modell w=2u l=2u
vd10 20 0 5
md10  21 19 0 0  modeld w=10u l=2u
ml10  20 20 21 0  modell w=2u l=2u
vd11 22 0 5
md11  23 21 0 0  modeld w=10u l=2u
ml11  22 22 23 0  modell w=2u l=2u
vd12 24 0 5
md12  25 23 0 0  modeld w=10u l=2u
ml12  24 24 25 0  modell w=2u l=2u
vd13 26 0 5
md13  27 25 0 0  modeld w=10u l=2u
ml13  26 26 27 0  modell w=2u l=2u
vd14 28 0 5
md14  29 27 0 0  modeld w=10u l=2u
ml14  28 28 29 0  modell w=2u l=2u
vd15 30 0 5
md15  31 29 0 0  modeld w=10u l=2u
ml15  30 30 31 0  modell w=2u l=2u
vd16 32 0 5
md16  33 31 0 0  modeld w=10u l=2u
ml16  32 32 33 0  modell w=2u l=2u
vd17 34 0 5
md17  35 33 0 0  modeld w=10u l=2u
ml17  34 34 35 0  modell w=2u l=2u
vd18 36 0 5
md18  37 35 0 0  modeld w=10u l=2u
ml18  36 36 37 0  modell w=2u l=2u
vd19 38 0 5
md19  39 37 0 0  modeld w=10u l=2u
ml19  38 38 39 0  modell w=2u l=2u
vd20 40 0 5
md20  41 39 0 0  modeld w=10u l=2u
ml20  40 40 41 0  modell w=2u l=2u
vd21 42 0 5
md21  43 41 0 0  modeld w=10u l=2u
ml21  42 42 43 0  modell w=2u l=2u
vd22 44 0 5
md22  45 43 0 0  modeld w=10u l=2u
ml22  44 44 45 0  modell w=2u l=2u
vd23 46 0 5
md23  47 45 0 0  modeld w=10u l=2u
ml23  46 46 47 0  modell w=2u l=2u
vd24 48 0 5
md24  49 47 0 0  modeld w=10u l=2u
ml24  48 48 49 0  modell w=2u l=2u
vd25 50 0 5
md25  51 49 0 0  modeld w=10u l=2u
ml25  50 50 51 0  modell w=2u l=2u
vd26 52 0 5
md26  53 51 0 0  modeld w=10u l=2u
ml26  52 52 53 0  modell w=2u l=2u
vd27 54 0 5
md27  55 53 0 0  modeld w=10u l=2u
ml27  54 54 55 0  modell w=2u l=2u
vd28 56 0 5
md28  57 55 0 0  modeld w=10u l=2u
ml28  56 56 57 0  modell w=2u l=2u
vd29 58 0 5
md29  59 57 0 0  modeld w=10u l=2u
ml29  58 58 59 0  modell w=2u l=2u
vd30 60 0 5
md30  61 59 0 0  modeld w=10u l=2u
ml30  60 60 61 0  modell w=2u l=2u
vd31 62 0 5
md31  63 61 0 0  modeld w=10u l=2u
ml31  62 62 63 0  modell w=2u l=2u
vd32 64 0 5
md32  65 63 0 0  modeld w=10u l=2u
ml32  64 64 65 0  modell w=2u l=2u
vd33 66 0 5
md33  67 65 0 0  modeld w=10u l=2u
ml33  66 66 67 0  modell w=2u l=2u
vd34 68 0 5
md34  69 67 0 0  modeld w=10u l=2u
ml34  68 68 69 0  modell w=2u l=2u
vd35 70 0 5
md35  71 69 0 0  modeld w=10u l=2u
ml35  70 70 71 0  modell w=2u l=2u
vd36 72 0 5
md36  73 71 0 0  modeld w=10u l=2u
ml36  72 72 73 0  modell w=2u l=2u
vd37 74 0 5
md37  75 73 0 0  modeld w=10u l=2u
ml37  74 74 75 0  modell w=2u l=2u
vd38 76 0 5
md38  77 75 0 0  modeld w=10u l=2u
ml38  76 76 77 0  modell w=2u l=2u
vd39 78 0 5
md39  79 77 0 0  modeld w=10u l=2u
ml39  78 78 79 0  modell w=2u l=2u
vd40 80 0 5
md40  81 79 0 0  modeld w=10u l=2u
ml40  80 80 81 0  modell w=2u l=2u
vd41 82 0 5
md41  83 81 0 0  modeld w=10u l=2u
ml41  82 82 83 0  modell w=2u l=2u
vd42 84 0 5
md42  85 83 0 0  modeld w=10u l=2u
ml42  84 84 85 0  modell w=2u l=2u
vd43 86 0 5
md43  87 85 0 0  modeld w=10u l=2u
ml43  86 86 87 0  modell w=2u l=2u
vd44 88 0 5
md44  89 87 0 0  modeld w=10u l=2u
ml44  88 88 89 0  modell w=2u l=2u
vd45 90 0 5
md45  91 89 0 0  modeld w=10u l=2u
ml45  90 90 91 0  modell w=2u l=2u
vd46 92 0 5
md46  93 91 0 0  modeld w=10u l=2u
ml46  92 92 93 0  modell w=2u l=2u
vd47 94 0 5
md47  95 93 0 0  modeld w=10u l=2u
ml47  94 94 95 0  modell w=2u l=2u
vd48 96 0 5
md48  97 95 0 0  modeld w=10u l=2u
ml48  96 96 97 0  modell w=2u l=2u
vd49 98 0 5
md49  99 97 0 0  modeld w=10u l=2u
ml49  98 98 99 0  modell w=2u l=2u
vd50 100 0 5
md50  101 99 0 0  modeld w=10u l=2u
ml50  100 100 101 0  modell w=2u l=2u
vd51 102 0 5
md51  103 101 0 0  modeld w=10u l=2u
ml51  102 102 103 0  modell w=2u l=2u
vd52 104 0 5
md52  105 103 0 0  modeld w=10u l=2u
ml52  104 104 105 0  modell w=2u l=2u
vd53 106 0 5
md53  107 105 0 0  modeld w=10u l=2u
ml53  106 106 107 0  modell w=2u l=2u
vd54 108 0 5
md54  109 107 0 0  modeld w=10u l=2u
ml54  108 108 109 0  modell w=2u l=2u
vd55 110 0 5
md55  111 109 0 0  modeld w=10u l=2u
ml55  110 110 111 0  modell w=2u l=2u
vd56 112 0 5
md56  113 111 0 0  modeld w=10u l=2u
ml56  112 112 113 0  modell w=2u l=2u
vd57 114 0 5
md57  115 113 0 0  modeld w=10u l=2u
ml57  114 114 115 0  modell w=2u l=2u
vd58 116 0 5
md58  117 115 0 0  modeld w=10u l=2u
ml58  116 116 117 0  modell w=2u l=2u
vd59 118 0 5
md59  119 117 0 0  modeld w=10u l=2u
ml59  118 118 119 0  modell w=2u l=2u
vd60 120 0 5
md60  121 119 0 0  modeld w=10u l=2u
ml60  120 120 121 0  modell w=2u l=2u
vd61 122 0 5
md61  123 121 0 0  modeld w=10u l=2u
ml61  122 122 123 0  modell w=2u l=2u
vd62 124 0 5
md62  125 123 0 0  modeld w=10u l=2u
ml62  124 124 125 0  modell w=2u l=2u
vd63 126 0 5
md63  127 125 0 0  modeld w=10u l=2u
ml63  126 126 127 0  modell w=2u l=2u
vd64 128 0 5
md64  129 127 0 0  modeld w=10u l=2u
ml64  128 128 129 0  modell w=2u l=2u
vd65 130 0 5
md65  131 129 0 0  modeld w=10u l=2u
ml65  130 130 131 0  modell w=2u l=2u
vd66 132 0 5
md66  133 131 0 0  modeld w=10u l=2u
ml66  132 132 133 0  modell w=2u l=2u
vd67 134 0 5
md67  135 133 0 0  modeld w=10u l=2u
ml67  134 134 135 0  modell w=2u l=2u
vd68 136 0 5
md68  137 135 0 0  modeld w=10u l=2u
ml68  136 136 137 0  modell w=2u l=2u
vd69 138 0 5
md69  139 137 0 0  modeld w=10u l=2u
ml69  138 138 139 0  modell w=2u l=2u
vd70 140 0 5
md70  141 139 0 0  modeld w=10u l=2u
ml70  140 140 141 0  modell w=2u l=2u
vd71 142 0 5
md71  143 141 0 0  modeld w=10u l=2u
ml71  142 142 143 0  modell w=2u l=2u
vd72 144 0 5
md72  145 143 0 0  modeld w=10u l=2u
ml72  144 144 145 0  modell w=2u l=2u
vd73 146 0 5
md73  147 145 0 0  modeld w=10u l=2u
ml73  146 146 147 0  modell w=2u l=2u
vd74 148 0 5
md74  149 147 0 0  modeld w=10u l=2u
ml74  148 148 149 0  modell w=2u l=2u
vd75 150 0 5
md75  151 149 0 0  modeld w=10u l=2u
ml75  150 150 151 0  modell w=2u l=2u
vd76 152 0 5
md76  153 151 0 0  modeld w=10u l=2u
ml76  152 152 153 0  modell w=2u l=2u
vd77 154 0 5
md77  155 153 0 0  modeld w=10u l=2u
ml77  154 154 155 0  modell w=2u l=2u
vd78 156 0 5
md78  157 155 0 0  modeld w=10u l=2u
ml78  156 156 157 0  modell w=2u l=2u
vd79 158 0 5
md79  159 157 0 0  modeld w=10u l=2u
ml79  158 158 159 0  modell w=2u l=2u
vd80 160 0 5
md80  161 159 0 0  modeld w=10u l=2u
ml80  160 160 161 0  modell w=2u l=2u
vd81 162 0 5
md81  163 161 0 0  modeld w=10u l=2u
ml81  162 162 163 0  modell w=2u l=2u
vd82 164 0 5
md82  165 163 0 0  modeld w=10u l=2u
ml82  164 164 165 0  modell w=2u l=2u
vd83 166 0 5
md83  167 165 0 0  modeld w=10u l=2u
ml83  166 166 167 0  modell w=2u l=2u
vd84 168 0 5
md84  169 167 0 0  modeld w=10u l=2u
ml84  168 168 169 0  modell w=2u l=2u
vd85 170 0 5
md85  171 169 0 0  modeld w=10u l=2u
ml85  170 170 171 0  modell w=2u l=2u
vd86 172 0 5
md86  173 171 0 0  modeld w=10u l=2u
ml86  172 172 173 0  modell w=2u l=2u
vd87 174 0 5
md87  175 173 0 0  modeld w=10u l=2u
ml87  174 174 175 0  modell w=2u l=2u
vd88 176 0 5
md88  177 175 0 0  modeld w=10u l=2u
ml88  176 176 177 0  modell w=2u l=2u
vd89 178 0 5
md89  179 177 0 0  modeld w=10u l=2u
ml89  178 178 179 0  modell w=2u l=2u
vd90 180 0 5
md90  181 179 0 0  modeld w=10u l=2u
ml90  180 180 181 0  modell w=2u l=2u
vd91 182 0 5
md91  183 181 0 0  modeld w=10u l=2u
ml91  182 182 183 0  modell w=2u l=2u
vd92 184 0 5
md92  185 183 0 0  modeld w=10u l=2u
ml92  184 184 185 0  modell w=2u l=2u
vd93 186 0 5
md93  187 185 0 0  modeld w=10u l=2u
ml93  186 186 187 0  modell w=2u l=2u
vd94 188 0 5
md94  189 187 0 0  modeld w=10u l=2u
ml94  188 188 189 0  modell w=2u l=2u
vd95 190 0 5
md95  191 189 0 0  modeld w=10u l=2u
ml95  190 190 191 0  modell w=2u l=2u
vd96 192 0 5
md96  193 191 0 0  modeld w=10u l=2u
ml96  192 192 193 0  modell w=2u l=2u
vd97 194 0 5
md97  195 193 0 0  modeld w=10u l=2u
ml97  194 194 195 0  modell w=2u l=2u
vd98 196 0 5
md98  197 195 0 0  modeld w=10u l=2u
ml98  196 196 197 0  modell w=2u l=2u
vd99 198 0 5
md99  199 197 0 0  modeld w=10u l=2u
ml99  198 198 199 0  modell w=2u l=2u
vd100 200 0 5
md100  201 199 0 0  modeld w=10u l=2u
ml100  200 200 201 0  modell w=2u l=2u
vin 1 0 .8
.MODEL MODELD NMOS (level=2 KP=28U VTO=0.7 LAMBDA=0.01 GAMMA=0.9 PHI=0.5)
.MODEL MODELL NMOS (level=2 KP=28U VTO=0.7 LAMBDA=0.01 GAMMA=0.9 PHI=0.5)
.width out=80
.PRINT OP iter(0) V(nodes)
.op
.end
