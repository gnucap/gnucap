Mutual inductance test circuit
v1 1 0  pulse(0 1 .002 .002 .002 .002 .01) ac 1
r1a 1 2 22
l1a 2 0 .56
l1b 3 0 .79
k1 l1a l1b .75
r1b 3 0 75

v2 4 0  pulse(0 1 .002 .002 .002 .002 .01) ac 1
r2a 4 5 22
l2a 5 6 .061151326
l2b 6 0 .498848674
l2c 6 7 .291151326
r2b 7 0 75

v3 8 0  pulse(0 1 .002 .002 .002 .002 .01) ac 1
r3a 8 9 22
l3a 10 0 .56
l3b 11 0 .79
e3a 9 10 11 0 .631454018
e3b 12 11 10 0 .890801204
r3b 12 0 75

.options nopage
.list
.width out=132
.print ac v(2) v(3) v(5) v(7) v(9) v(12)
.ac dec 2 .1 1k
.print tran v(2) v(3) v(5) v(7) v(9) v(12)
.tran .001 .01 0 .0001
.list
.status notime
.end
