'
v1 1 0 1
e1 2 0 1 0  pwl(-5 -2 -3 0 0 0 4 1)
e2 3 0 1 0  pwl(-5 -2 -3 0 -3 1 0 0 4 1)
e3 4 0 1 0  pwl(-5 -2 -3 0 0 -3 4 5)
'e4 5 0 1 0  pwl(4 1 0 0 -3 0 -5 2)
.option out=170
.print dc v(nodes) f(e*) ev(e*)
.dc v1 -10 10 .5
.end
