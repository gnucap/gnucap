# voltage source test
v1 0 1 1 ac 1
r1 1 2 1k
r2 0 2 1k
e1 0 3 0 2 4.
r3 0 3 1k
g1 0 4 0 2 4.
r3 0 4 1k
.list
.print op v(1) v(2) v(3) v(4)
.op
.print op vo(e1) vin(e1) i(e1) p(e1) pd(e1) ps(e1)
.op
.print op vo(v1) vin(v1) i(v1) p(v1) pd(v1) ps(v1)
.op
.print ac v(1) v(2) v(3) v(4)
.ac 1k
.print ac vo(e1) vin(e1) i(e1) p(e1) pd(e1) ps(e1)
.ac 1k
.print ac vo(v1) vin(v1) i(v1) p(v1) pd(v1) ps(v1)
.ac 1k
.end
