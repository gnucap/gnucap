;'trunc error check
V1   1  0  ac 1 pwl (0 0 1p 1)
L3   1  2  .1
R4   2  0  1.
R5   1  3  1.
C6   3  0  .1
.options short=1p trtol=7 reltol=.01 method=euler
.width out=170
.list
.print tran iter(0)  v(nodes) z(c6) zraw(c6) z(3) control(0) timef(C6) timef(L3) dt(C6) dtr(C6)
.tran 0 .1 .01 trace rejected
* exact=0.632120559
.list
.status notime
.end
