'6 inverters as gates
.gen freq=1 offset=2.5 init=2.5 ampl=2.5 
Vdd  8  0  dc 5.
V1   1  0  generator( 1. ) 
U2   2 0 8 8 1  mos inv
U3   3 0 8 8 2  mos inv
U4   4 0 8 8 3  mos inv
U5   5 0 8 8 4  mos inv
U6   6 0 8 8 5  mos inv
U7   7 0 8 8 6  mos inv
.model  mos logic ( delay= 1n  rise= 1n  fall= 1n  rs= 100.  rw= 1.G 
+ thh= 0.75  thl= 0.25  mr= 5.  mf= 5.  over=10k vmax= 5.  vmin= 0. )
.subckt mosinv1  2  4  1  5  3 
M1   2  3  4  4  nmos  l= 100.u  w= 100.u  nrd= 1.  nrs= 1. 
M2   2  3  1  1  pmos  l= 100.u  w= 100.u  nrd= 1.  nrs= 1. 
.ends
*+ends mosinv1
.model nmos  nmos ( level=2  vto= 0.  gamma= 0.  phi= 0.6  is= 10.E-15 pb= 0.8 
+ cgso= 0.  cgdo= 0.  cgbo= 0.  rsh= 0.  cj= 0.  mj= 0.5  cjsw= 0.  mjsw= 0.33 
+ tox= 100.n  nfs= 0.  tpg=1  ld= 0.  uo= 600.  neff= 1.  fc= 0.5  delta= 0. 
+)
*+(* vfb=-0.6 * kp= 20.71886u )
.model pmos  pmos ( level=2  vto= 0.  gamma= 0.  phi= 0.6  is= 10.E-15 pb= 0.8 
+ cgso= 0.  cgdo= 0.  cgbo= 0.  rsh= 0.  cj= 0.  mj= 0.5  cjsw= 0.  mjsw= 0.33 
+ tox= 100.n  nfs= 0.  tpg=1  ld= 0.  uo= 600.  neff= 1.  fc= 0.5  delta= 0. 
+)
*+(* vfb=-0.6 * kp= 20.71886u )
.option mode=mixed vmax=5.1 vmin=-.1
.print op v(1 2 3 4 5 6 7 8) logic(1 2 3 4 5 6 7 8)
.op
'.option trace
'.print tran v(nodes) l(nodes)
'.tran 0 10 .05 
.stat notime
.end 
