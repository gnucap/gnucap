# coil errors
l1 1 0 1
r2 2 0 1
k1 l1 r2 .9
.print ac v(nodes)
.ac 1k
.end
