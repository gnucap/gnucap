' exp test
.option out=170
.param delay=10n
v1 1 0 exp  iv= 0.  pv= 1.  td1=delay/10  tau1=delay/2  td2=delay  tau2=delay/2
.print tran v 1
.tran 0 'delay*2' 'delay/200'
.list
.end
