'trunc error check
V1   1  0  generator(1)
L3   1  2  .1
R4   2  0  1.
R5   1  3  1.
C6   3  0  .1
.options short=1p trtol=7 reltol=.001
.width out=170
.list
.print tran iter(0)  v(nodes) i(L3) i(R4) control(0)
.fanout
.fanout 2
.tran 0 .1 .01 trace rejected
.print ac v(nodes) vp(nodes) i(L3) i(R4) ip(L3) ip(R4) -v(1) vp(1)
.ac .001 100 decade 2
.list
.status notime
.end
