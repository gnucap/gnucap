100 cascaded NMOS inverters
md1  3 2 0 0  modeld w=10u l=2u
ml1  1 1 3 0  modell w=2u l=2u
md2  4 3 0 0  modeld w=10u l=2u
ml2  1 1 4 0  modell w=2u l=2u
md3  5 4 0 0  modeld w=10u l=2u
ml3  1 1 5 0  modell w=2u l=2u
md4  6 5 0 0  modeld w=10u l=2u
ml4  1 1 6 0  modell w=2u l=2u
md5  7 6 0 0  modeld w=10u l=2u
ml5  1 1 7 0  modell w=2u l=2u
md6  8 7 0 0  modeld w=10u l=2u
ml6  1 1 8 0  modell w=2u l=2u
md7  9 8 0 0  modeld w=10u l=2u
ml7  1 1 9 0  modell w=2u l=2u
md8  10 9 0 0  modeld w=10u l=2u
ml8  1 1 10 0  modell w=2u l=2u
md9  11 10 0 0  modeld w=10u l=2u
ml9  1 1 11 0  modell w=2u l=2u
md10  12 11 0 0  modeld w=10u l=2u
ml10  1 1 12 0  modell w=2u l=2u
md11  13 12 0 0  modeld w=10u l=2u
ml11  1 1 13 0  modell w=2u l=2u
md12  14 13 0 0  modeld w=10u l=2u
ml12  1 1 14 0  modell w=2u l=2u
md13  15 14 0 0  modeld w=10u l=2u
ml13  1 1 15 0  modell w=2u l=2u
md14  16 15 0 0  modeld w=10u l=2u
ml14  1 1 16 0  modell w=2u l=2u
md15  17 16 0 0  modeld w=10u l=2u
ml15  1 1 17 0  modell w=2u l=2u
md16  18 17 0 0  modeld w=10u l=2u
ml16  1 1 18 0  modell w=2u l=2u
md17  19 18 0 0  modeld w=10u l=2u
ml17  1 1 19 0  modell w=2u l=2u
md18  20 19 0 0  modeld w=10u l=2u
ml18  1 1 20 0  modell w=2u l=2u
md19  21 20 0 0  modeld w=10u l=2u
ml19  1 1 21 0  modell w=2u l=2u
md20  22 21 0 0  modeld w=10u l=2u
ml20  1 1 22 0  modell w=2u l=2u
md21  23 22 0 0  modeld w=10u l=2u
ml21  1 1 23 0  modell w=2u l=2u
md22  24 23 0 0  modeld w=10u l=2u
ml22  1 1 24 0  modell w=2u l=2u
md23  25 24 0 0  modeld w=10u l=2u
ml23  1 1 25 0  modell w=2u l=2u
md24  26 25 0 0  modeld w=10u l=2u
ml24  1 1 26 0  modell w=2u l=2u
md25  27 26 0 0  modeld w=10u l=2u
ml25  1 1 27 0  modell w=2u l=2u
md26  28 27 0 0  modeld w=10u l=2u
ml26  1 1 28 0  modell w=2u l=2u
md27  29 28 0 0  modeld w=10u l=2u
ml27  1 1 29 0  modell w=2u l=2u
md28  30 29 0 0  modeld w=10u l=2u
ml28  1 1 30 0  modell w=2u l=2u
md29  31 30 0 0  modeld w=10u l=2u
ml29  1 1 31 0  modell w=2u l=2u
md30  32 31 0 0  modeld w=10u l=2u
ml30  1 1 32 0  modell w=2u l=2u
md31  33 32 0 0  modeld w=10u l=2u
ml31  1 1 33 0  modell w=2u l=2u
md32  34 33 0 0  modeld w=10u l=2u
ml32  1 1 34 0  modell w=2u l=2u
md33  35 34 0 0  modeld w=10u l=2u
ml33  1 1 35 0  modell w=2u l=2u
md34  36 35 0 0  modeld w=10u l=2u
ml34  1 1 36 0  modell w=2u l=2u
md35  37 36 0 0  modeld w=10u l=2u
ml35  1 1 37 0  modell w=2u l=2u
md36  38 37 0 0  modeld w=10u l=2u
ml36  1 1 38 0  modell w=2u l=2u
md37  39 38 0 0  modeld w=10u l=2u
ml37  1 1 39 0  modell w=2u l=2u
md38  40 39 0 0  modeld w=10u l=2u
ml38  1 1 40 0  modell w=2u l=2u
md39  41 40 0 0  modeld w=10u l=2u
ml39  1 1 41 0  modell w=2u l=2u
md40  42 41 0 0  modeld w=10u l=2u
ml40  1 1 42 0  modell w=2u l=2u
md41  43 42 0 0  modeld w=10u l=2u
ml41  1 1 43 0  modell w=2u l=2u
md42  44 43 0 0  modeld w=10u l=2u
ml42  1 1 44 0  modell w=2u l=2u
md43  45 44 0 0  modeld w=10u l=2u
ml43  1 1 45 0  modell w=2u l=2u
md44  46 45 0 0  modeld w=10u l=2u
ml44  1 1 46 0  modell w=2u l=2u
md45  47 46 0 0  modeld w=10u l=2u
ml45  1 1 47 0  modell w=2u l=2u
md46  48 47 0 0  modeld w=10u l=2u
ml46  1 1 48 0  modell w=2u l=2u
md47  49 48 0 0  modeld w=10u l=2u
ml47  1 1 49 0  modell w=2u l=2u
md48  50 49 0 0  modeld w=10u l=2u
ml48  1 1 50 0  modell w=2u l=2u
md49  51 50 0 0  modeld w=10u l=2u
ml49  1 1 51 0  modell w=2u l=2u
md50  52 51 0 0  modeld w=10u l=2u
ml50  1 1 52 0  modell w=2u l=2u
md51  53 52 0 0  modeld w=10u l=2u
ml51  1 1 53 0  modell w=2u l=2u
md52  54 53 0 0  modeld w=10u l=2u
ml52  1 1 54 0  modell w=2u l=2u
md53  55 54 0 0  modeld w=10u l=2u
ml53  1 1 55 0  modell w=2u l=2u
md54  56 55 0 0  modeld w=10u l=2u
ml54  1 1 56 0  modell w=2u l=2u
md55  57 56 0 0  modeld w=10u l=2u
ml55  1 1 57 0  modell w=2u l=2u
md56  58 57 0 0  modeld w=10u l=2u
ml56  1 1 58 0  modell w=2u l=2u
md57  59 58 0 0  modeld w=10u l=2u
ml57  1 1 59 0  modell w=2u l=2u
md58  60 59 0 0  modeld w=10u l=2u
ml58  1 1 60 0  modell w=2u l=2u
md59  61 60 0 0  modeld w=10u l=2u
ml59  1 1 61 0  modell w=2u l=2u
md60  62 61 0 0  modeld w=10u l=2u
ml60  1 1 62 0  modell w=2u l=2u
md61  63 62 0 0  modeld w=10u l=2u
ml61  1 1 63 0  modell w=2u l=2u
md62  64 63 0 0  modeld w=10u l=2u
ml62  1 1 64 0  modell w=2u l=2u
md63  65 64 0 0  modeld w=10u l=2u
ml63  1 1 65 0  modell w=2u l=2u
md64  66 65 0 0  modeld w=10u l=2u
ml64  1 1 66 0  modell w=2u l=2u
md65  67 66 0 0  modeld w=10u l=2u
ml65  1 1 67 0  modell w=2u l=2u
md66  68 67 0 0  modeld w=10u l=2u
ml66  1 1 68 0  modell w=2u l=2u
md67  69 68 0 0  modeld w=10u l=2u
ml67  1 1 69 0  modell w=2u l=2u
md68  70 69 0 0  modeld w=10u l=2u
ml68  1 1 70 0  modell w=2u l=2u
md69  71 70 0 0  modeld w=10u l=2u
ml69  1 1 71 0  modell w=2u l=2u
md70  72 71 0 0  modeld w=10u l=2u
ml70  1 1 72 0  modell w=2u l=2u
md71  73 72 0 0  modeld w=10u l=2u
ml71  1 1 73 0  modell w=2u l=2u
md72  74 73 0 0  modeld w=10u l=2u
ml72  1 1 74 0  modell w=2u l=2u
md73  75 74 0 0  modeld w=10u l=2u
ml73  1 1 75 0  modell w=2u l=2u
md74  76 75 0 0  modeld w=10u l=2u
ml74  1 1 76 0  modell w=2u l=2u
md75  77 76 0 0  modeld w=10u l=2u
ml75  1 1 77 0  modell w=2u l=2u
md76  78 77 0 0  modeld w=10u l=2u
ml76  1 1 78 0  modell w=2u l=2u
md77  79 78 0 0  modeld w=10u l=2u
ml77  1 1 79 0  modell w=2u l=2u
md78  80 79 0 0  modeld w=10u l=2u
ml78  1 1 80 0  modell w=2u l=2u
md79  81 80 0 0  modeld w=10u l=2u
ml79  1 1 81 0  modell w=2u l=2u
md80  82 81 0 0  modeld w=10u l=2u
ml80  1 1 82 0  modell w=2u l=2u
md81  83 82 0 0  modeld w=10u l=2u
ml81  1 1 83 0  modell w=2u l=2u
md82  84 83 0 0  modeld w=10u l=2u
ml82  1 1 84 0  modell w=2u l=2u
md83  85 84 0 0  modeld w=10u l=2u
ml83  1 1 85 0  modell w=2u l=2u
md84  86 85 0 0  modeld w=10u l=2u
ml84  1 1 86 0  modell w=2u l=2u
md85  87 86 0 0  modeld w=10u l=2u
ml85  1 1 87 0  modell w=2u l=2u
md86  88 87 0 0  modeld w=10u l=2u
ml86  1 1 88 0  modell w=2u l=2u
md87  89 88 0 0  modeld w=10u l=2u
ml87  1 1 89 0  modell w=2u l=2u
md88  90 89 0 0  modeld w=10u l=2u
ml88  1 1 90 0  modell w=2u l=2u
md89  91 90 0 0  modeld w=10u l=2u
ml89  1 1 91 0  modell w=2u l=2u
md90  92 91 0 0  modeld w=10u l=2u
ml90  1 1 92 0  modell w=2u l=2u
md91  93 92 0 0  modeld w=10u l=2u
ml91  1 1 93 0  modell w=2u l=2u
md92  94 93 0 0  modeld w=10u l=2u
ml92  1 1 94 0  modell w=2u l=2u
md93  95 94 0 0  modeld w=10u l=2u
ml93  1 1 95 0  modell w=2u l=2u
md94  96 95 0 0  modeld w=10u l=2u
ml94  1 1 96 0  modell w=2u l=2u
md95  97 96 0 0  modeld w=10u l=2u
ml95  1 1 97 0  modell w=2u l=2u
md96  98 97 0 0  modeld w=10u l=2u
ml96  1 1 98 0  modell w=2u l=2u
md97  99 98 0 0  modeld w=10u l=2u
ml97  1 1 99 0  modell w=2u l=2u
md98  100 99 0 0  modeld w=10u l=2u
ml98  1 1 100 0  modell w=2u l=2u
md99  101 100 0 0  modeld w=10u l=2u
ml99  1 1 101 0  modell w=2u l=2u
md100  102 101 0 0  modeld w=10u l=2u
ml100  1 1 102 0  modell w=2u l=2u
vdd 1 0 5
vin 2 0 .8
.MODEL MODELD NMOS (level=2 KP=28U VTO=0.7 LAMBDA=0.01 GAMMA=0.9 PHI=0.5)
.MODEL MODELL NMOS (level=2 KP=28U VTO=0.7 LAMBDA=0.01 GAMMA=0.9 PHI=0.5)
.width out=80
.PRINT OP iter(0) V(nodes)
.option vmin=-.1 short=1u dampstrategy=10
.op
.end
