30x30 grid test

.subckt grids top1 top900 bot450
.parameter r=1
.parameter l=1e-6
.parameter c=1e-9
Rtop_1_2 top1 top2 {r}
Ltop_1_2 top1 top2 {l}
Rbot_1_2 bot1 bot2 {r}
Lbot_1_2 bot1 bot2 {l}
Rtop_1_31 top1 top31 {r}
Ltop_1_31 top1 top31 {l}
Rbot_1_31 bot1 bot31 {r}
Lbot_1_31 bot1 bot31 {l}
C1 top1 bot1 {c}
Rtop_2_3 top2 top3 {r}
Ltop_2_3 top2 top3 {l}
Rbot_2_3 bot2 bot3 {r}
Lbot_2_3 bot2 bot3 {l}
Rtop_2_32 top2 top32 {r}
Ltop_2_32 top2 top32 {l}
Rbot_2_32 bot2 bot32 {r}
Lbot_2_32 bot2 bot32 {l}
C2 top2 bot2 {c}
Rtop_3_4 top3 top4 {r}
Ltop_3_4 top3 top4 {l}
Rbot_3_4 bot3 bot4 {r}
Lbot_3_4 bot3 bot4 {l}
Rtop_3_33 top3 top33 {r}
Ltop_3_33 top3 top33 {l}
Rbot_3_33 bot3 bot33 {r}
Lbot_3_33 bot3 bot33 {l}
C3 top3 bot3 {c}
Rtop_4_5 top4 top5 {r}
Ltop_4_5 top4 top5 {l}
Rbot_4_5 bot4 bot5 {r}
Lbot_4_5 bot4 bot5 {l}
Rtop_4_34 top4 top34 {r}
Ltop_4_34 top4 top34 {l}
Rbot_4_34 bot4 bot34 {r}
Lbot_4_34 bot4 bot34 {l}
C4 top4 bot4 {c}
Rtop_5_6 top5 top6 {r}
Ltop_5_6 top5 top6 {l}
Rbot_5_6 bot5 bot6 {r}
Lbot_5_6 bot5 bot6 {l}
Rtop_5_35 top5 top35 {r}
Ltop_5_35 top5 top35 {l}
Rbot_5_35 bot5 bot35 {r}
Lbot_5_35 bot5 bot35 {l}
C5 top5 bot5 {c}
Rtop_6_7 top6 top7 {r}
Ltop_6_7 top6 top7 {l}
Rbot_6_7 bot6 bot7 {r}
Lbot_6_7 bot6 bot7 {l}
Rtop_6_36 top6 top36 {r}
Ltop_6_36 top6 top36 {l}
Rbot_6_36 bot6 bot36 {r}
Lbot_6_36 bot6 bot36 {l}
C6 top6 bot6 {c}
Rtop_7_8 top7 top8 {r}
Ltop_7_8 top7 top8 {l}
Rbot_7_8 bot7 bot8 {r}
Lbot_7_8 bot7 bot8 {l}
Rtop_7_37 top7 top37 {r}
Ltop_7_37 top7 top37 {l}
Rbot_7_37 bot7 bot37 {r}
Lbot_7_37 bot7 bot37 {l}
C7 top7 bot7 {c}
Rtop_8_9 top8 top9 {r}
Ltop_8_9 top8 top9 {l}
Rbot_8_9 bot8 bot9 {r}
Lbot_8_9 bot8 bot9 {l}
Rtop_8_38 top8 top38 {r}
Ltop_8_38 top8 top38 {l}
Rbot_8_38 bot8 bot38 {r}
Lbot_8_38 bot8 bot38 {l}
C8 top8 bot8 {c}
Rtop_9_10 top9 top10 {r}
Ltop_9_10 top9 top10 {l}
Rbot_9_10 bot9 bot10 {r}
Lbot_9_10 bot9 bot10 {l}
Rtop_9_39 top9 top39 {r}
Ltop_9_39 top9 top39 {l}
Rbot_9_39 bot9 bot39 {r}
Lbot_9_39 bot9 bot39 {l}
C9 top9 bot9 {c}
Rtop_10_11 top10 top11 {r}
Ltop_10_11 top10 top11 {l}
Rbot_10_11 bot10 bot11 {r}
Lbot_10_11 bot10 bot11 {l}
Rtop_10_40 top10 top40 {r}
Ltop_10_40 top10 top40 {l}
Rbot_10_40 bot10 bot40 {r}
Lbot_10_40 bot10 bot40 {l}
C10 top10 bot10 {c}
Rtop_11_12 top11 top12 {r}
Ltop_11_12 top11 top12 {l}
Rbot_11_12 bot11 bot12 {r}
Lbot_11_12 bot11 bot12 {l}
Rtop_11_41 top11 top41 {r}
Ltop_11_41 top11 top41 {l}
Rbot_11_41 bot11 bot41 {r}
Lbot_11_41 bot11 bot41 {l}
C11 top11 bot11 {c}
Rtop_12_13 top12 top13 {r}
Ltop_12_13 top12 top13 {l}
Rbot_12_13 bot12 bot13 {r}
Lbot_12_13 bot12 bot13 {l}
Rtop_12_42 top12 top42 {r}
Ltop_12_42 top12 top42 {l}
Rbot_12_42 bot12 bot42 {r}
Lbot_12_42 bot12 bot42 {l}
C12 top12 bot12 {c}
Rtop_13_14 top13 top14 {r}
Ltop_13_14 top13 top14 {l}
Rbot_13_14 bot13 bot14 {r}
Lbot_13_14 bot13 bot14 {l}
Rtop_13_43 top13 top43 {r}
Ltop_13_43 top13 top43 {l}
Rbot_13_43 bot13 bot43 {r}
Lbot_13_43 bot13 bot43 {l}
C13 top13 bot13 {c}
Rtop_14_15 top14 top15 {r}
Ltop_14_15 top14 top15 {l}
Rbot_14_15 bot14 bot15 {r}
Lbot_14_15 bot14 bot15 {l}
Rtop_14_44 top14 top44 {r}
Ltop_14_44 top14 top44 {l}
Rbot_14_44 bot14 bot44 {r}
Lbot_14_44 bot14 bot44 {l}
C14 top14 bot14 {c}
Rtop_15_16 top15 top16 {r}
Ltop_15_16 top15 top16 {l}
Rbot_15_16 bot15 bot16 {r}
Lbot_15_16 bot15 bot16 {l}
Rtop_15_45 top15 top45 {r}
Ltop_15_45 top15 top45 {l}
Rbot_15_45 bot15 bot45 {r}
Lbot_15_45 bot15 bot45 {l}
C15 top15 bot15 {c}
Rtop_16_17 top16 top17 {r}
Ltop_16_17 top16 top17 {l}
Rbot_16_17 bot16 bot17 {r}
Lbot_16_17 bot16 bot17 {l}
Rtop_16_46 top16 top46 {r}
Ltop_16_46 top16 top46 {l}
Rbot_16_46 bot16 bot46 {r}
Lbot_16_46 bot16 bot46 {l}
C16 top16 bot16 {c}
Rtop_17_18 top17 top18 {r}
Ltop_17_18 top17 top18 {l}
Rbot_17_18 bot17 bot18 {r}
Lbot_17_18 bot17 bot18 {l}
Rtop_17_47 top17 top47 {r}
Ltop_17_47 top17 top47 {l}
Rbot_17_47 bot17 bot47 {r}
Lbot_17_47 bot17 bot47 {l}
C17 top17 bot17 {c}
Rtop_18_19 top18 top19 {r}
Ltop_18_19 top18 top19 {l}
Rbot_18_19 bot18 bot19 {r}
Lbot_18_19 bot18 bot19 {l}
Rtop_18_48 top18 top48 {r}
Ltop_18_48 top18 top48 {l}
Rbot_18_48 bot18 bot48 {r}
Lbot_18_48 bot18 bot48 {l}
C18 top18 bot18 {c}
Rtop_19_20 top19 top20 {r}
Ltop_19_20 top19 top20 {l}
Rbot_19_20 bot19 bot20 {r}
Lbot_19_20 bot19 bot20 {l}
Rtop_19_49 top19 top49 {r}
Ltop_19_49 top19 top49 {l}
Rbot_19_49 bot19 bot49 {r}
Lbot_19_49 bot19 bot49 {l}
C19 top19 bot19 {c}
Rtop_20_21 top20 top21 {r}
Ltop_20_21 top20 top21 {l}
Rbot_20_21 bot20 bot21 {r}
Lbot_20_21 bot20 bot21 {l}
Rtop_20_50 top20 top50 {r}
Ltop_20_50 top20 top50 {l}
Rbot_20_50 bot20 bot50 {r}
Lbot_20_50 bot20 bot50 {l}
C20 top20 bot20 {c}
Rtop_21_22 top21 top22 {r}
Ltop_21_22 top21 top22 {l}
Rbot_21_22 bot21 bot22 {r}
Lbot_21_22 bot21 bot22 {l}
Rtop_21_51 top21 top51 {r}
Ltop_21_51 top21 top51 {l}
Rbot_21_51 bot21 bot51 {r}
Lbot_21_51 bot21 bot51 {l}
C21 top21 bot21 {c}
Rtop_22_23 top22 top23 {r}
Ltop_22_23 top22 top23 {l}
Rbot_22_23 bot22 bot23 {r}
Lbot_22_23 bot22 bot23 {l}
Rtop_22_52 top22 top52 {r}
Ltop_22_52 top22 top52 {l}
Rbot_22_52 bot22 bot52 {r}
Lbot_22_52 bot22 bot52 {l}
C22 top22 bot22 {c}
Rtop_23_24 top23 top24 {r}
Ltop_23_24 top23 top24 {l}
Rbot_23_24 bot23 bot24 {r}
Lbot_23_24 bot23 bot24 {l}
Rtop_23_53 top23 top53 {r}
Ltop_23_53 top23 top53 {l}
Rbot_23_53 bot23 bot53 {r}
Lbot_23_53 bot23 bot53 {l}
C23 top23 bot23 {c}
Rtop_24_25 top24 top25 {r}
Ltop_24_25 top24 top25 {l}
Rbot_24_25 bot24 bot25 {r}
Lbot_24_25 bot24 bot25 {l}
Rtop_24_54 top24 top54 {r}
Ltop_24_54 top24 top54 {l}
Rbot_24_54 bot24 bot54 {r}
Lbot_24_54 bot24 bot54 {l}
C24 top24 bot24 {c}
Rtop_25_26 top25 top26 {r}
Ltop_25_26 top25 top26 {l}
Rbot_25_26 bot25 bot26 {r}
Lbot_25_26 bot25 bot26 {l}
Rtop_25_55 top25 top55 {r}
Ltop_25_55 top25 top55 {l}
Rbot_25_55 bot25 bot55 {r}
Lbot_25_55 bot25 bot55 {l}
C25 top25 bot25 {c}
Rtop_26_27 top26 top27 {r}
Ltop_26_27 top26 top27 {l}
Rbot_26_27 bot26 bot27 {r}
Lbot_26_27 bot26 bot27 {l}
Rtop_26_56 top26 top56 {r}
Ltop_26_56 top26 top56 {l}
Rbot_26_56 bot26 bot56 {r}
Lbot_26_56 bot26 bot56 {l}
C26 top26 bot26 {c}
Rtop_27_28 top27 top28 {r}
Ltop_27_28 top27 top28 {l}
Rbot_27_28 bot27 bot28 {r}
Lbot_27_28 bot27 bot28 {l}
Rtop_27_57 top27 top57 {r}
Ltop_27_57 top27 top57 {l}
Rbot_27_57 bot27 bot57 {r}
Lbot_27_57 bot27 bot57 {l}
C27 top27 bot27 {c}
Rtop_28_29 top28 top29 {r}
Ltop_28_29 top28 top29 {l}
Rbot_28_29 bot28 bot29 {r}
Lbot_28_29 bot28 bot29 {l}
Rtop_28_58 top28 top58 {r}
Ltop_28_58 top28 top58 {l}
Rbot_28_58 bot28 bot58 {r}
Lbot_28_58 bot28 bot58 {l}
C28 top28 bot28 {c}
Rtop_29_30 top29 top30 {r}
Ltop_29_30 top29 top30 {l}
Rbot_29_30 bot29 bot30 {r}
Lbot_29_30 bot29 bot30 {l}
Rtop_29_59 top29 top59 {r}
Ltop_29_59 top29 top59 {l}
Rbot_29_59 bot29 bot59 {r}
Lbot_29_59 bot29 bot59 {l}
C29 top29 bot29 {c}
Rtop_30_60 top30 top60 {r}
Ltop_30_60 top30 top60 {l}
Rbot_30_60 bot30 bot60 {r}
Lbot_30_60 bot30 bot60 {l}
C30 top30 bot30 {c}
Rtop_31_32 top31 top32 {r}
Ltop_31_32 top31 top32 {l}
Rbot_31_32 bot31 bot32 {r}
Lbot_31_32 bot31 bot32 {l}
Rtop_31_61 top31 top61 {r}
Ltop_31_61 top31 top61 {l}
Rbot_31_61 bot31 bot61 {r}
Lbot_31_61 bot31 bot61 {l}
C31 top31 bot31 {c}
Rtop_32_33 top32 top33 {r}
Ltop_32_33 top32 top33 {l}
Rbot_32_33 bot32 bot33 {r}
Lbot_32_33 bot32 bot33 {l}
Rtop_32_62 top32 top62 {r}
Ltop_32_62 top32 top62 {l}
Rbot_32_62 bot32 bot62 {r}
Lbot_32_62 bot32 bot62 {l}
C32 top32 bot32 {c}
Rtop_33_34 top33 top34 {r}
Ltop_33_34 top33 top34 {l}
Rbot_33_34 bot33 bot34 {r}
Lbot_33_34 bot33 bot34 {l}
Rtop_33_63 top33 top63 {r}
Ltop_33_63 top33 top63 {l}
Rbot_33_63 bot33 bot63 {r}
Lbot_33_63 bot33 bot63 {l}
C33 top33 bot33 {c}
Rtop_34_35 top34 top35 {r}
Ltop_34_35 top34 top35 {l}
Rbot_34_35 bot34 bot35 {r}
Lbot_34_35 bot34 bot35 {l}
Rtop_34_64 top34 top64 {r}
Ltop_34_64 top34 top64 {l}
Rbot_34_64 bot34 bot64 {r}
Lbot_34_64 bot34 bot64 {l}
C34 top34 bot34 {c}
Rtop_35_36 top35 top36 {r}
Ltop_35_36 top35 top36 {l}
Rbot_35_36 bot35 bot36 {r}
Lbot_35_36 bot35 bot36 {l}
Rtop_35_65 top35 top65 {r}
Ltop_35_65 top35 top65 {l}
Rbot_35_65 bot35 bot65 {r}
Lbot_35_65 bot35 bot65 {l}
C35 top35 bot35 {c}
Rtop_36_37 top36 top37 {r}
Ltop_36_37 top36 top37 {l}
Rbot_36_37 bot36 bot37 {r}
Lbot_36_37 bot36 bot37 {l}
Rtop_36_66 top36 top66 {r}
Ltop_36_66 top36 top66 {l}
Rbot_36_66 bot36 bot66 {r}
Lbot_36_66 bot36 bot66 {l}
C36 top36 bot36 {c}
Rtop_37_38 top37 top38 {r}
Ltop_37_38 top37 top38 {l}
Rbot_37_38 bot37 bot38 {r}
Lbot_37_38 bot37 bot38 {l}
Rtop_37_67 top37 top67 {r}
Ltop_37_67 top37 top67 {l}
Rbot_37_67 bot37 bot67 {r}
Lbot_37_67 bot37 bot67 {l}
C37 top37 bot37 {c}
Rtop_38_39 top38 top39 {r}
Ltop_38_39 top38 top39 {l}
Rbot_38_39 bot38 bot39 {r}
Lbot_38_39 bot38 bot39 {l}
Rtop_38_68 top38 top68 {r}
Ltop_38_68 top38 top68 {l}
Rbot_38_68 bot38 bot68 {r}
Lbot_38_68 bot38 bot68 {l}
C38 top38 bot38 {c}
Rtop_39_40 top39 top40 {r}
Ltop_39_40 top39 top40 {l}
Rbot_39_40 bot39 bot40 {r}
Lbot_39_40 bot39 bot40 {l}
Rtop_39_69 top39 top69 {r}
Ltop_39_69 top39 top69 {l}
Rbot_39_69 bot39 bot69 {r}
Lbot_39_69 bot39 bot69 {l}
C39 top39 bot39 {c}
Rtop_40_41 top40 top41 {r}
Ltop_40_41 top40 top41 {l}
Rbot_40_41 bot40 bot41 {r}
Lbot_40_41 bot40 bot41 {l}
Rtop_40_70 top40 top70 {r}
Ltop_40_70 top40 top70 {l}
Rbot_40_70 bot40 bot70 {r}
Lbot_40_70 bot40 bot70 {l}
C40 top40 bot40 {c}
Rtop_41_42 top41 top42 {r}
Ltop_41_42 top41 top42 {l}
Rbot_41_42 bot41 bot42 {r}
Lbot_41_42 bot41 bot42 {l}
Rtop_41_71 top41 top71 {r}
Ltop_41_71 top41 top71 {l}
Rbot_41_71 bot41 bot71 {r}
Lbot_41_71 bot41 bot71 {l}
C41 top41 bot41 {c}
Rtop_42_43 top42 top43 {r}
Ltop_42_43 top42 top43 {l}
Rbot_42_43 bot42 bot43 {r}
Lbot_42_43 bot42 bot43 {l}
Rtop_42_72 top42 top72 {r}
Ltop_42_72 top42 top72 {l}
Rbot_42_72 bot42 bot72 {r}
Lbot_42_72 bot42 bot72 {l}
C42 top42 bot42 {c}
Rtop_43_44 top43 top44 {r}
Ltop_43_44 top43 top44 {l}
Rbot_43_44 bot43 bot44 {r}
Lbot_43_44 bot43 bot44 {l}
Rtop_43_73 top43 top73 {r}
Ltop_43_73 top43 top73 {l}
Rbot_43_73 bot43 bot73 {r}
Lbot_43_73 bot43 bot73 {l}
C43 top43 bot43 {c}
Rtop_44_45 top44 top45 {r}
Ltop_44_45 top44 top45 {l}
Rbot_44_45 bot44 bot45 {r}
Lbot_44_45 bot44 bot45 {l}
Rtop_44_74 top44 top74 {r}
Ltop_44_74 top44 top74 {l}
Rbot_44_74 bot44 bot74 {r}
Lbot_44_74 bot44 bot74 {l}
C44 top44 bot44 {c}
Rtop_45_46 top45 top46 {r}
Ltop_45_46 top45 top46 {l}
Rbot_45_46 bot45 bot46 {r}
Lbot_45_46 bot45 bot46 {l}
Rtop_45_75 top45 top75 {r}
Ltop_45_75 top45 top75 {l}
Rbot_45_75 bot45 bot75 {r}
Lbot_45_75 bot45 bot75 {l}
C45 top45 bot45 {c}
Rtop_46_47 top46 top47 {r}
Ltop_46_47 top46 top47 {l}
Rbot_46_47 bot46 bot47 {r}
Lbot_46_47 bot46 bot47 {l}
Rtop_46_76 top46 top76 {r}
Ltop_46_76 top46 top76 {l}
Rbot_46_76 bot46 bot76 {r}
Lbot_46_76 bot46 bot76 {l}
C46 top46 bot46 {c}
Rtop_47_48 top47 top48 {r}
Ltop_47_48 top47 top48 {l}
Rbot_47_48 bot47 bot48 {r}
Lbot_47_48 bot47 bot48 {l}
Rtop_47_77 top47 top77 {r}
Ltop_47_77 top47 top77 {l}
Rbot_47_77 bot47 bot77 {r}
Lbot_47_77 bot47 bot77 {l}
C47 top47 bot47 {c}
Rtop_48_49 top48 top49 {r}
Ltop_48_49 top48 top49 {l}
Rbot_48_49 bot48 bot49 {r}
Lbot_48_49 bot48 bot49 {l}
Rtop_48_78 top48 top78 {r}
Ltop_48_78 top48 top78 {l}
Rbot_48_78 bot48 bot78 {r}
Lbot_48_78 bot48 bot78 {l}
C48 top48 bot48 {c}
Rtop_49_50 top49 top50 {r}
Ltop_49_50 top49 top50 {l}
Rbot_49_50 bot49 bot50 {r}
Lbot_49_50 bot49 bot50 {l}
Rtop_49_79 top49 top79 {r}
Ltop_49_79 top49 top79 {l}
Rbot_49_79 bot49 bot79 {r}
Lbot_49_79 bot49 bot79 {l}
C49 top49 bot49 {c}
Rtop_50_51 top50 top51 {r}
Ltop_50_51 top50 top51 {l}
Rbot_50_51 bot50 bot51 {r}
Lbot_50_51 bot50 bot51 {l}
Rtop_50_80 top50 top80 {r}
Ltop_50_80 top50 top80 {l}
Rbot_50_80 bot50 bot80 {r}
Lbot_50_80 bot50 bot80 {l}
C50 top50 bot50 {c}
Rtop_51_52 top51 top52 {r}
Ltop_51_52 top51 top52 {l}
Rbot_51_52 bot51 bot52 {r}
Lbot_51_52 bot51 bot52 {l}
Rtop_51_81 top51 top81 {r}
Ltop_51_81 top51 top81 {l}
Rbot_51_81 bot51 bot81 {r}
Lbot_51_81 bot51 bot81 {l}
C51 top51 bot51 {c}
Rtop_52_53 top52 top53 {r}
Ltop_52_53 top52 top53 {l}
Rbot_52_53 bot52 bot53 {r}
Lbot_52_53 bot52 bot53 {l}
Rtop_52_82 top52 top82 {r}
Ltop_52_82 top52 top82 {l}
Rbot_52_82 bot52 bot82 {r}
Lbot_52_82 bot52 bot82 {l}
C52 top52 bot52 {c}
Rtop_53_54 top53 top54 {r}
Ltop_53_54 top53 top54 {l}
Rbot_53_54 bot53 bot54 {r}
Lbot_53_54 bot53 bot54 {l}
Rtop_53_83 top53 top83 {r}
Ltop_53_83 top53 top83 {l}
Rbot_53_83 bot53 bot83 {r}
Lbot_53_83 bot53 bot83 {l}
C53 top53 bot53 {c}
Rtop_54_55 top54 top55 {r}
Ltop_54_55 top54 top55 {l}
Rbot_54_55 bot54 bot55 {r}
Lbot_54_55 bot54 bot55 {l}
Rtop_54_84 top54 top84 {r}
Ltop_54_84 top54 top84 {l}
Rbot_54_84 bot54 bot84 {r}
Lbot_54_84 bot54 bot84 {l}
C54 top54 bot54 {c}
Rtop_55_56 top55 top56 {r}
Ltop_55_56 top55 top56 {l}
Rbot_55_56 bot55 bot56 {r}
Lbot_55_56 bot55 bot56 {l}
Rtop_55_85 top55 top85 {r}
Ltop_55_85 top55 top85 {l}
Rbot_55_85 bot55 bot85 {r}
Lbot_55_85 bot55 bot85 {l}
C55 top55 bot55 {c}
Rtop_56_57 top56 top57 {r}
Ltop_56_57 top56 top57 {l}
Rbot_56_57 bot56 bot57 {r}
Lbot_56_57 bot56 bot57 {l}
Rtop_56_86 top56 top86 {r}
Ltop_56_86 top56 top86 {l}
Rbot_56_86 bot56 bot86 {r}
Lbot_56_86 bot56 bot86 {l}
C56 top56 bot56 {c}
Rtop_57_58 top57 top58 {r}
Ltop_57_58 top57 top58 {l}
Rbot_57_58 bot57 bot58 {r}
Lbot_57_58 bot57 bot58 {l}
Rtop_57_87 top57 top87 {r}
Ltop_57_87 top57 top87 {l}
Rbot_57_87 bot57 bot87 {r}
Lbot_57_87 bot57 bot87 {l}
C57 top57 bot57 {c}
Rtop_58_59 top58 top59 {r}
Ltop_58_59 top58 top59 {l}
Rbot_58_59 bot58 bot59 {r}
Lbot_58_59 bot58 bot59 {l}
Rtop_58_88 top58 top88 {r}
Ltop_58_88 top58 top88 {l}
Rbot_58_88 bot58 bot88 {r}
Lbot_58_88 bot58 bot88 {l}
C58 top58 bot58 {c}
Rtop_59_60 top59 top60 {r}
Ltop_59_60 top59 top60 {l}
Rbot_59_60 bot59 bot60 {r}
Lbot_59_60 bot59 bot60 {l}
Rtop_59_89 top59 top89 {r}
Ltop_59_89 top59 top89 {l}
Rbot_59_89 bot59 bot89 {r}
Lbot_59_89 bot59 bot89 {l}
C59 top59 bot59 {c}
Rtop_60_90 top60 top90 {r}
Ltop_60_90 top60 top90 {l}
Rbot_60_90 bot60 bot90 {r}
Lbot_60_90 bot60 bot90 {l}
C60 top60 bot60 {c}
Rtop_61_62 top61 top62 {r}
Ltop_61_62 top61 top62 {l}
Rbot_61_62 bot61 bot62 {r}
Lbot_61_62 bot61 bot62 {l}
Rtop_61_91 top61 top91 {r}
Ltop_61_91 top61 top91 {l}
Rbot_61_91 bot61 bot91 {r}
Lbot_61_91 bot61 bot91 {l}
C61 top61 bot61 {c}
Rtop_62_63 top62 top63 {r}
Ltop_62_63 top62 top63 {l}
Rbot_62_63 bot62 bot63 {r}
Lbot_62_63 bot62 bot63 {l}
Rtop_62_92 top62 top92 {r}
Ltop_62_92 top62 top92 {l}
Rbot_62_92 bot62 bot92 {r}
Lbot_62_92 bot62 bot92 {l}
C62 top62 bot62 {c}
Rtop_63_64 top63 top64 {r}
Ltop_63_64 top63 top64 {l}
Rbot_63_64 bot63 bot64 {r}
Lbot_63_64 bot63 bot64 {l}
Rtop_63_93 top63 top93 {r}
Ltop_63_93 top63 top93 {l}
Rbot_63_93 bot63 bot93 {r}
Lbot_63_93 bot63 bot93 {l}
C63 top63 bot63 {c}
Rtop_64_65 top64 top65 {r}
Ltop_64_65 top64 top65 {l}
Rbot_64_65 bot64 bot65 {r}
Lbot_64_65 bot64 bot65 {l}
Rtop_64_94 top64 top94 {r}
Ltop_64_94 top64 top94 {l}
Rbot_64_94 bot64 bot94 {r}
Lbot_64_94 bot64 bot94 {l}
C64 top64 bot64 {c}
Rtop_65_66 top65 top66 {r}
Ltop_65_66 top65 top66 {l}
Rbot_65_66 bot65 bot66 {r}
Lbot_65_66 bot65 bot66 {l}
Rtop_65_95 top65 top95 {r}
Ltop_65_95 top65 top95 {l}
Rbot_65_95 bot65 bot95 {r}
Lbot_65_95 bot65 bot95 {l}
C65 top65 bot65 {c}
Rtop_66_67 top66 top67 {r}
Ltop_66_67 top66 top67 {l}
Rbot_66_67 bot66 bot67 {r}
Lbot_66_67 bot66 bot67 {l}
Rtop_66_96 top66 top96 {r}
Ltop_66_96 top66 top96 {l}
Rbot_66_96 bot66 bot96 {r}
Lbot_66_96 bot66 bot96 {l}
C66 top66 bot66 {c}
Rtop_67_68 top67 top68 {r}
Ltop_67_68 top67 top68 {l}
Rbot_67_68 bot67 bot68 {r}
Lbot_67_68 bot67 bot68 {l}
Rtop_67_97 top67 top97 {r}
Ltop_67_97 top67 top97 {l}
Rbot_67_97 bot67 bot97 {r}
Lbot_67_97 bot67 bot97 {l}
C67 top67 bot67 {c}
Rtop_68_69 top68 top69 {r}
Ltop_68_69 top68 top69 {l}
Rbot_68_69 bot68 bot69 {r}
Lbot_68_69 bot68 bot69 {l}
Rtop_68_98 top68 top98 {r}
Ltop_68_98 top68 top98 {l}
Rbot_68_98 bot68 bot98 {r}
Lbot_68_98 bot68 bot98 {l}
C68 top68 bot68 {c}
Rtop_69_70 top69 top70 {r}
Ltop_69_70 top69 top70 {l}
Rbot_69_70 bot69 bot70 {r}
Lbot_69_70 bot69 bot70 {l}
Rtop_69_99 top69 top99 {r}
Ltop_69_99 top69 top99 {l}
Rbot_69_99 bot69 bot99 {r}
Lbot_69_99 bot69 bot99 {l}
C69 top69 bot69 {c}
Rtop_70_71 top70 top71 {r}
Ltop_70_71 top70 top71 {l}
Rbot_70_71 bot70 bot71 {r}
Lbot_70_71 bot70 bot71 {l}
Rtop_70_100 top70 top100 {r}
Ltop_70_100 top70 top100 {l}
Rbot_70_100 bot70 bot100 {r}
Lbot_70_100 bot70 bot100 {l}
C70 top70 bot70 {c}
Rtop_71_72 top71 top72 {r}
Ltop_71_72 top71 top72 {l}
Rbot_71_72 bot71 bot72 {r}
Lbot_71_72 bot71 bot72 {l}
Rtop_71_101 top71 top101 {r}
Ltop_71_101 top71 top101 {l}
Rbot_71_101 bot71 bot101 {r}
Lbot_71_101 bot71 bot101 {l}
C71 top71 bot71 {c}
Rtop_72_73 top72 top73 {r}
Ltop_72_73 top72 top73 {l}
Rbot_72_73 bot72 bot73 {r}
Lbot_72_73 bot72 bot73 {l}
Rtop_72_102 top72 top102 {r}
Ltop_72_102 top72 top102 {l}
Rbot_72_102 bot72 bot102 {r}
Lbot_72_102 bot72 bot102 {l}
C72 top72 bot72 {c}
Rtop_73_74 top73 top74 {r}
Ltop_73_74 top73 top74 {l}
Rbot_73_74 bot73 bot74 {r}
Lbot_73_74 bot73 bot74 {l}
Rtop_73_103 top73 top103 {r}
Ltop_73_103 top73 top103 {l}
Rbot_73_103 bot73 bot103 {r}
Lbot_73_103 bot73 bot103 {l}
C73 top73 bot73 {c}
Rtop_74_75 top74 top75 {r}
Ltop_74_75 top74 top75 {l}
Rbot_74_75 bot74 bot75 {r}
Lbot_74_75 bot74 bot75 {l}
Rtop_74_104 top74 top104 {r}
Ltop_74_104 top74 top104 {l}
Rbot_74_104 bot74 bot104 {r}
Lbot_74_104 bot74 bot104 {l}
C74 top74 bot74 {c}
Rtop_75_76 top75 top76 {r}
Ltop_75_76 top75 top76 {l}
Rbot_75_76 bot75 bot76 {r}
Lbot_75_76 bot75 bot76 {l}
Rtop_75_105 top75 top105 {r}
Ltop_75_105 top75 top105 {l}
Rbot_75_105 bot75 bot105 {r}
Lbot_75_105 bot75 bot105 {l}
C75 top75 bot75 {c}
Rtop_76_77 top76 top77 {r}
Ltop_76_77 top76 top77 {l}
Rbot_76_77 bot76 bot77 {r}
Lbot_76_77 bot76 bot77 {l}
Rtop_76_106 top76 top106 {r}
Ltop_76_106 top76 top106 {l}
Rbot_76_106 bot76 bot106 {r}
Lbot_76_106 bot76 bot106 {l}
C76 top76 bot76 {c}
Rtop_77_78 top77 top78 {r}
Ltop_77_78 top77 top78 {l}
Rbot_77_78 bot77 bot78 {r}
Lbot_77_78 bot77 bot78 {l}
Rtop_77_107 top77 top107 {r}
Ltop_77_107 top77 top107 {l}
Rbot_77_107 bot77 bot107 {r}
Lbot_77_107 bot77 bot107 {l}
C77 top77 bot77 {c}
Rtop_78_79 top78 top79 {r}
Ltop_78_79 top78 top79 {l}
Rbot_78_79 bot78 bot79 {r}
Lbot_78_79 bot78 bot79 {l}
Rtop_78_108 top78 top108 {r}
Ltop_78_108 top78 top108 {l}
Rbot_78_108 bot78 bot108 {r}
Lbot_78_108 bot78 bot108 {l}
C78 top78 bot78 {c}
Rtop_79_80 top79 top80 {r}
Ltop_79_80 top79 top80 {l}
Rbot_79_80 bot79 bot80 {r}
Lbot_79_80 bot79 bot80 {l}
Rtop_79_109 top79 top109 {r}
Ltop_79_109 top79 top109 {l}
Rbot_79_109 bot79 bot109 {r}
Lbot_79_109 bot79 bot109 {l}
C79 top79 bot79 {c}
Rtop_80_81 top80 top81 {r}
Ltop_80_81 top80 top81 {l}
Rbot_80_81 bot80 bot81 {r}
Lbot_80_81 bot80 bot81 {l}
Rtop_80_110 top80 top110 {r}
Ltop_80_110 top80 top110 {l}
Rbot_80_110 bot80 bot110 {r}
Lbot_80_110 bot80 bot110 {l}
C80 top80 bot80 {c}
Rtop_81_82 top81 top82 {r}
Ltop_81_82 top81 top82 {l}
Rbot_81_82 bot81 bot82 {r}
Lbot_81_82 bot81 bot82 {l}
Rtop_81_111 top81 top111 {r}
Ltop_81_111 top81 top111 {l}
Rbot_81_111 bot81 bot111 {r}
Lbot_81_111 bot81 bot111 {l}
C81 top81 bot81 {c}
Rtop_82_83 top82 top83 {r}
Ltop_82_83 top82 top83 {l}
Rbot_82_83 bot82 bot83 {r}
Lbot_82_83 bot82 bot83 {l}
Rtop_82_112 top82 top112 {r}
Ltop_82_112 top82 top112 {l}
Rbot_82_112 bot82 bot112 {r}
Lbot_82_112 bot82 bot112 {l}
C82 top82 bot82 {c}
Rtop_83_84 top83 top84 {r}
Ltop_83_84 top83 top84 {l}
Rbot_83_84 bot83 bot84 {r}
Lbot_83_84 bot83 bot84 {l}
Rtop_83_113 top83 top113 {r}
Ltop_83_113 top83 top113 {l}
Rbot_83_113 bot83 bot113 {r}
Lbot_83_113 bot83 bot113 {l}
C83 top83 bot83 {c}
Rtop_84_85 top84 top85 {r}
Ltop_84_85 top84 top85 {l}
Rbot_84_85 bot84 bot85 {r}
Lbot_84_85 bot84 bot85 {l}
Rtop_84_114 top84 top114 {r}
Ltop_84_114 top84 top114 {l}
Rbot_84_114 bot84 bot114 {r}
Lbot_84_114 bot84 bot114 {l}
C84 top84 bot84 {c}
Rtop_85_86 top85 top86 {r}
Ltop_85_86 top85 top86 {l}
Rbot_85_86 bot85 bot86 {r}
Lbot_85_86 bot85 bot86 {l}
Rtop_85_115 top85 top115 {r}
Ltop_85_115 top85 top115 {l}
Rbot_85_115 bot85 bot115 {r}
Lbot_85_115 bot85 bot115 {l}
C85 top85 bot85 {c}
Rtop_86_87 top86 top87 {r}
Ltop_86_87 top86 top87 {l}
Rbot_86_87 bot86 bot87 {r}
Lbot_86_87 bot86 bot87 {l}
Rtop_86_116 top86 top116 {r}
Ltop_86_116 top86 top116 {l}
Rbot_86_116 bot86 bot116 {r}
Lbot_86_116 bot86 bot116 {l}
C86 top86 bot86 {c}
Rtop_87_88 top87 top88 {r}
Ltop_87_88 top87 top88 {l}
Rbot_87_88 bot87 bot88 {r}
Lbot_87_88 bot87 bot88 {l}
Rtop_87_117 top87 top117 {r}
Ltop_87_117 top87 top117 {l}
Rbot_87_117 bot87 bot117 {r}
Lbot_87_117 bot87 bot117 {l}
C87 top87 bot87 {c}
Rtop_88_89 top88 top89 {r}
Ltop_88_89 top88 top89 {l}
Rbot_88_89 bot88 bot89 {r}
Lbot_88_89 bot88 bot89 {l}
Rtop_88_118 top88 top118 {r}
Ltop_88_118 top88 top118 {l}
Rbot_88_118 bot88 bot118 {r}
Lbot_88_118 bot88 bot118 {l}
C88 top88 bot88 {c}
Rtop_89_90 top89 top90 {r}
Ltop_89_90 top89 top90 {l}
Rbot_89_90 bot89 bot90 {r}
Lbot_89_90 bot89 bot90 {l}
Rtop_89_119 top89 top119 {r}
Ltop_89_119 top89 top119 {l}
Rbot_89_119 bot89 bot119 {r}
Lbot_89_119 bot89 bot119 {l}
C89 top89 bot89 {c}
Rtop_90_120 top90 top120 {r}
Ltop_90_120 top90 top120 {l}
Rbot_90_120 bot90 bot120 {r}
Lbot_90_120 bot90 bot120 {l}
C90 top90 bot90 {c}
Rtop_91_92 top91 top92 {r}
Ltop_91_92 top91 top92 {l}
Rbot_91_92 bot91 bot92 {r}
Lbot_91_92 bot91 bot92 {l}
Rtop_91_121 top91 top121 {r}
Ltop_91_121 top91 top121 {l}
Rbot_91_121 bot91 bot121 {r}
Lbot_91_121 bot91 bot121 {l}
C91 top91 bot91 {c}
Rtop_92_93 top92 top93 {r}
Ltop_92_93 top92 top93 {l}
Rbot_92_93 bot92 bot93 {r}
Lbot_92_93 bot92 bot93 {l}
Rtop_92_122 top92 top122 {r}
Ltop_92_122 top92 top122 {l}
Rbot_92_122 bot92 bot122 {r}
Lbot_92_122 bot92 bot122 {l}
C92 top92 bot92 {c}
Rtop_93_94 top93 top94 {r}
Ltop_93_94 top93 top94 {l}
Rbot_93_94 bot93 bot94 {r}
Lbot_93_94 bot93 bot94 {l}
Rtop_93_123 top93 top123 {r}
Ltop_93_123 top93 top123 {l}
Rbot_93_123 bot93 bot123 {r}
Lbot_93_123 bot93 bot123 {l}
C93 top93 bot93 {c}
Rtop_94_95 top94 top95 {r}
Ltop_94_95 top94 top95 {l}
Rbot_94_95 bot94 bot95 {r}
Lbot_94_95 bot94 bot95 {l}
Rtop_94_124 top94 top124 {r}
Ltop_94_124 top94 top124 {l}
Rbot_94_124 bot94 bot124 {r}
Lbot_94_124 bot94 bot124 {l}
C94 top94 bot94 {c}
Rtop_95_96 top95 top96 {r}
Ltop_95_96 top95 top96 {l}
Rbot_95_96 bot95 bot96 {r}
Lbot_95_96 bot95 bot96 {l}
Rtop_95_125 top95 top125 {r}
Ltop_95_125 top95 top125 {l}
Rbot_95_125 bot95 bot125 {r}
Lbot_95_125 bot95 bot125 {l}
C95 top95 bot95 {c}
Rtop_96_97 top96 top97 {r}
Ltop_96_97 top96 top97 {l}
Rbot_96_97 bot96 bot97 {r}
Lbot_96_97 bot96 bot97 {l}
Rtop_96_126 top96 top126 {r}
Ltop_96_126 top96 top126 {l}
Rbot_96_126 bot96 bot126 {r}
Lbot_96_126 bot96 bot126 {l}
C96 top96 bot96 {c}
Rtop_97_98 top97 top98 {r}
Ltop_97_98 top97 top98 {l}
Rbot_97_98 bot97 bot98 {r}
Lbot_97_98 bot97 bot98 {l}
Rtop_97_127 top97 top127 {r}
Ltop_97_127 top97 top127 {l}
Rbot_97_127 bot97 bot127 {r}
Lbot_97_127 bot97 bot127 {l}
C97 top97 bot97 {c}
Rtop_98_99 top98 top99 {r}
Ltop_98_99 top98 top99 {l}
Rbot_98_99 bot98 bot99 {r}
Lbot_98_99 bot98 bot99 {l}
Rtop_98_128 top98 top128 {r}
Ltop_98_128 top98 top128 {l}
Rbot_98_128 bot98 bot128 {r}
Lbot_98_128 bot98 bot128 {l}
C98 top98 bot98 {c}
Rtop_99_100 top99 top100 {r}
Ltop_99_100 top99 top100 {l}
Rbot_99_100 bot99 bot100 {r}
Lbot_99_100 bot99 bot100 {l}
Rtop_99_129 top99 top129 {r}
Ltop_99_129 top99 top129 {l}
Rbot_99_129 bot99 bot129 {r}
Lbot_99_129 bot99 bot129 {l}
C99 top99 bot99 {c}
Rtop_100_101 top100 top101 {r}
Ltop_100_101 top100 top101 {l}
Rbot_100_101 bot100 bot101 {r}
Lbot_100_101 bot100 bot101 {l}
Rtop_100_130 top100 top130 {r}
Ltop_100_130 top100 top130 {l}
Rbot_100_130 bot100 bot130 {r}
Lbot_100_130 bot100 bot130 {l}
C100 top100 bot100 {c}
Rtop_101_102 top101 top102 {r}
Ltop_101_102 top101 top102 {l}
Rbot_101_102 bot101 bot102 {r}
Lbot_101_102 bot101 bot102 {l}
Rtop_101_131 top101 top131 {r}
Ltop_101_131 top101 top131 {l}
Rbot_101_131 bot101 bot131 {r}
Lbot_101_131 bot101 bot131 {l}
C101 top101 bot101 {c}
Rtop_102_103 top102 top103 {r}
Ltop_102_103 top102 top103 {l}
Rbot_102_103 bot102 bot103 {r}
Lbot_102_103 bot102 bot103 {l}
Rtop_102_132 top102 top132 {r}
Ltop_102_132 top102 top132 {l}
Rbot_102_132 bot102 bot132 {r}
Lbot_102_132 bot102 bot132 {l}
C102 top102 bot102 {c}
Rtop_103_104 top103 top104 {r}
Ltop_103_104 top103 top104 {l}
Rbot_103_104 bot103 bot104 {r}
Lbot_103_104 bot103 bot104 {l}
Rtop_103_133 top103 top133 {r}
Ltop_103_133 top103 top133 {l}
Rbot_103_133 bot103 bot133 {r}
Lbot_103_133 bot103 bot133 {l}
C103 top103 bot103 {c}
Rtop_104_105 top104 top105 {r}
Ltop_104_105 top104 top105 {l}
Rbot_104_105 bot104 bot105 {r}
Lbot_104_105 bot104 bot105 {l}
Rtop_104_134 top104 top134 {r}
Ltop_104_134 top104 top134 {l}
Rbot_104_134 bot104 bot134 {r}
Lbot_104_134 bot104 bot134 {l}
C104 top104 bot104 {c}
Rtop_105_106 top105 top106 {r}
Ltop_105_106 top105 top106 {l}
Rbot_105_106 bot105 bot106 {r}
Lbot_105_106 bot105 bot106 {l}
Rtop_105_135 top105 top135 {r}
Ltop_105_135 top105 top135 {l}
Rbot_105_135 bot105 bot135 {r}
Lbot_105_135 bot105 bot135 {l}
C105 top105 bot105 {c}
Rtop_106_107 top106 top107 {r}
Ltop_106_107 top106 top107 {l}
Rbot_106_107 bot106 bot107 {r}
Lbot_106_107 bot106 bot107 {l}
Rtop_106_136 top106 top136 {r}
Ltop_106_136 top106 top136 {l}
Rbot_106_136 bot106 bot136 {r}
Lbot_106_136 bot106 bot136 {l}
C106 top106 bot106 {c}
Rtop_107_108 top107 top108 {r}
Ltop_107_108 top107 top108 {l}
Rbot_107_108 bot107 bot108 {r}
Lbot_107_108 bot107 bot108 {l}
Rtop_107_137 top107 top137 {r}
Ltop_107_137 top107 top137 {l}
Rbot_107_137 bot107 bot137 {r}
Lbot_107_137 bot107 bot137 {l}
C107 top107 bot107 {c}
Rtop_108_109 top108 top109 {r}
Ltop_108_109 top108 top109 {l}
Rbot_108_109 bot108 bot109 {r}
Lbot_108_109 bot108 bot109 {l}
Rtop_108_138 top108 top138 {r}
Ltop_108_138 top108 top138 {l}
Rbot_108_138 bot108 bot138 {r}
Lbot_108_138 bot108 bot138 {l}
C108 top108 bot108 {c}
Rtop_109_110 top109 top110 {r}
Ltop_109_110 top109 top110 {l}
Rbot_109_110 bot109 bot110 {r}
Lbot_109_110 bot109 bot110 {l}
Rtop_109_139 top109 top139 {r}
Ltop_109_139 top109 top139 {l}
Rbot_109_139 bot109 bot139 {r}
Lbot_109_139 bot109 bot139 {l}
C109 top109 bot109 {c}
Rtop_110_111 top110 top111 {r}
Ltop_110_111 top110 top111 {l}
Rbot_110_111 bot110 bot111 {r}
Lbot_110_111 bot110 bot111 {l}
Rtop_110_140 top110 top140 {r}
Ltop_110_140 top110 top140 {l}
Rbot_110_140 bot110 bot140 {r}
Lbot_110_140 bot110 bot140 {l}
C110 top110 bot110 {c}
Rtop_111_112 top111 top112 {r}
Ltop_111_112 top111 top112 {l}
Rbot_111_112 bot111 bot112 {r}
Lbot_111_112 bot111 bot112 {l}
Rtop_111_141 top111 top141 {r}
Ltop_111_141 top111 top141 {l}
Rbot_111_141 bot111 bot141 {r}
Lbot_111_141 bot111 bot141 {l}
C111 top111 bot111 {c}
Rtop_112_113 top112 top113 {r}
Ltop_112_113 top112 top113 {l}
Rbot_112_113 bot112 bot113 {r}
Lbot_112_113 bot112 bot113 {l}
Rtop_112_142 top112 top142 {r}
Ltop_112_142 top112 top142 {l}
Rbot_112_142 bot112 bot142 {r}
Lbot_112_142 bot112 bot142 {l}
C112 top112 bot112 {c}
Rtop_113_114 top113 top114 {r}
Ltop_113_114 top113 top114 {l}
Rbot_113_114 bot113 bot114 {r}
Lbot_113_114 bot113 bot114 {l}
Rtop_113_143 top113 top143 {r}
Ltop_113_143 top113 top143 {l}
Rbot_113_143 bot113 bot143 {r}
Lbot_113_143 bot113 bot143 {l}
C113 top113 bot113 {c}
Rtop_114_115 top114 top115 {r}
Ltop_114_115 top114 top115 {l}
Rbot_114_115 bot114 bot115 {r}
Lbot_114_115 bot114 bot115 {l}
Rtop_114_144 top114 top144 {r}
Ltop_114_144 top114 top144 {l}
Rbot_114_144 bot114 bot144 {r}
Lbot_114_144 bot114 bot144 {l}
C114 top114 bot114 {c}
Rtop_115_116 top115 top116 {r}
Ltop_115_116 top115 top116 {l}
Rbot_115_116 bot115 bot116 {r}
Lbot_115_116 bot115 bot116 {l}
Rtop_115_145 top115 top145 {r}
Ltop_115_145 top115 top145 {l}
Rbot_115_145 bot115 bot145 {r}
Lbot_115_145 bot115 bot145 {l}
C115 top115 bot115 {c}
Rtop_116_117 top116 top117 {r}
Ltop_116_117 top116 top117 {l}
Rbot_116_117 bot116 bot117 {r}
Lbot_116_117 bot116 bot117 {l}
Rtop_116_146 top116 top146 {r}
Ltop_116_146 top116 top146 {l}
Rbot_116_146 bot116 bot146 {r}
Lbot_116_146 bot116 bot146 {l}
C116 top116 bot116 {c}
Rtop_117_118 top117 top118 {r}
Ltop_117_118 top117 top118 {l}
Rbot_117_118 bot117 bot118 {r}
Lbot_117_118 bot117 bot118 {l}
Rtop_117_147 top117 top147 {r}
Ltop_117_147 top117 top147 {l}
Rbot_117_147 bot117 bot147 {r}
Lbot_117_147 bot117 bot147 {l}
C117 top117 bot117 {c}
Rtop_118_119 top118 top119 {r}
Ltop_118_119 top118 top119 {l}
Rbot_118_119 bot118 bot119 {r}
Lbot_118_119 bot118 bot119 {l}
Rtop_118_148 top118 top148 {r}
Ltop_118_148 top118 top148 {l}
Rbot_118_148 bot118 bot148 {r}
Lbot_118_148 bot118 bot148 {l}
C118 top118 bot118 {c}
Rtop_119_120 top119 top120 {r}
Ltop_119_120 top119 top120 {l}
Rbot_119_120 bot119 bot120 {r}
Lbot_119_120 bot119 bot120 {l}
Rtop_119_149 top119 top149 {r}
Ltop_119_149 top119 top149 {l}
Rbot_119_149 bot119 bot149 {r}
Lbot_119_149 bot119 bot149 {l}
C119 top119 bot119 {c}
Rtop_120_150 top120 top150 {r}
Ltop_120_150 top120 top150 {l}
Rbot_120_150 bot120 bot150 {r}
Lbot_120_150 bot120 bot150 {l}
C120 top120 bot120 {c}
Rtop_121_122 top121 top122 {r}
Ltop_121_122 top121 top122 {l}
Rbot_121_122 bot121 bot122 {r}
Lbot_121_122 bot121 bot122 {l}
Rtop_121_151 top121 top151 {r}
Ltop_121_151 top121 top151 {l}
Rbot_121_151 bot121 bot151 {r}
Lbot_121_151 bot121 bot151 {l}
C121 top121 bot121 {c}
Rtop_122_123 top122 top123 {r}
Ltop_122_123 top122 top123 {l}
Rbot_122_123 bot122 bot123 {r}
Lbot_122_123 bot122 bot123 {l}
Rtop_122_152 top122 top152 {r}
Ltop_122_152 top122 top152 {l}
Rbot_122_152 bot122 bot152 {r}
Lbot_122_152 bot122 bot152 {l}
C122 top122 bot122 {c}
Rtop_123_124 top123 top124 {r}
Ltop_123_124 top123 top124 {l}
Rbot_123_124 bot123 bot124 {r}
Lbot_123_124 bot123 bot124 {l}
Rtop_123_153 top123 top153 {r}
Ltop_123_153 top123 top153 {l}
Rbot_123_153 bot123 bot153 {r}
Lbot_123_153 bot123 bot153 {l}
C123 top123 bot123 {c}
Rtop_124_125 top124 top125 {r}
Ltop_124_125 top124 top125 {l}
Rbot_124_125 bot124 bot125 {r}
Lbot_124_125 bot124 bot125 {l}
Rtop_124_154 top124 top154 {r}
Ltop_124_154 top124 top154 {l}
Rbot_124_154 bot124 bot154 {r}
Lbot_124_154 bot124 bot154 {l}
C124 top124 bot124 {c}
Rtop_125_126 top125 top126 {r}
Ltop_125_126 top125 top126 {l}
Rbot_125_126 bot125 bot126 {r}
Lbot_125_126 bot125 bot126 {l}
Rtop_125_155 top125 top155 {r}
Ltop_125_155 top125 top155 {l}
Rbot_125_155 bot125 bot155 {r}
Lbot_125_155 bot125 bot155 {l}
C125 top125 bot125 {c}
Rtop_126_127 top126 top127 {r}
Ltop_126_127 top126 top127 {l}
Rbot_126_127 bot126 bot127 {r}
Lbot_126_127 bot126 bot127 {l}
Rtop_126_156 top126 top156 {r}
Ltop_126_156 top126 top156 {l}
Rbot_126_156 bot126 bot156 {r}
Lbot_126_156 bot126 bot156 {l}
C126 top126 bot126 {c}
Rtop_127_128 top127 top128 {r}
Ltop_127_128 top127 top128 {l}
Rbot_127_128 bot127 bot128 {r}
Lbot_127_128 bot127 bot128 {l}
Rtop_127_157 top127 top157 {r}
Ltop_127_157 top127 top157 {l}
Rbot_127_157 bot127 bot157 {r}
Lbot_127_157 bot127 bot157 {l}
C127 top127 bot127 {c}
Rtop_128_129 top128 top129 {r}
Ltop_128_129 top128 top129 {l}
Rbot_128_129 bot128 bot129 {r}
Lbot_128_129 bot128 bot129 {l}
Rtop_128_158 top128 top158 {r}
Ltop_128_158 top128 top158 {l}
Rbot_128_158 bot128 bot158 {r}
Lbot_128_158 bot128 bot158 {l}
C128 top128 bot128 {c}
Rtop_129_130 top129 top130 {r}
Ltop_129_130 top129 top130 {l}
Rbot_129_130 bot129 bot130 {r}
Lbot_129_130 bot129 bot130 {l}
Rtop_129_159 top129 top159 {r}
Ltop_129_159 top129 top159 {l}
Rbot_129_159 bot129 bot159 {r}
Lbot_129_159 bot129 bot159 {l}
C129 top129 bot129 {c}
Rtop_130_131 top130 top131 {r}
Ltop_130_131 top130 top131 {l}
Rbot_130_131 bot130 bot131 {r}
Lbot_130_131 bot130 bot131 {l}
Rtop_130_160 top130 top160 {r}
Ltop_130_160 top130 top160 {l}
Rbot_130_160 bot130 bot160 {r}
Lbot_130_160 bot130 bot160 {l}
C130 top130 bot130 {c}
Rtop_131_132 top131 top132 {r}
Ltop_131_132 top131 top132 {l}
Rbot_131_132 bot131 bot132 {r}
Lbot_131_132 bot131 bot132 {l}
Rtop_131_161 top131 top161 {r}
Ltop_131_161 top131 top161 {l}
Rbot_131_161 bot131 bot161 {r}
Lbot_131_161 bot131 bot161 {l}
C131 top131 bot131 {c}
Rtop_132_133 top132 top133 {r}
Ltop_132_133 top132 top133 {l}
Rbot_132_133 bot132 bot133 {r}
Lbot_132_133 bot132 bot133 {l}
Rtop_132_162 top132 top162 {r}
Ltop_132_162 top132 top162 {l}
Rbot_132_162 bot132 bot162 {r}
Lbot_132_162 bot132 bot162 {l}
C132 top132 bot132 {c}
Rtop_133_134 top133 top134 {r}
Ltop_133_134 top133 top134 {l}
Rbot_133_134 bot133 bot134 {r}
Lbot_133_134 bot133 bot134 {l}
Rtop_133_163 top133 top163 {r}
Ltop_133_163 top133 top163 {l}
Rbot_133_163 bot133 bot163 {r}
Lbot_133_163 bot133 bot163 {l}
C133 top133 bot133 {c}
Rtop_134_135 top134 top135 {r}
Ltop_134_135 top134 top135 {l}
Rbot_134_135 bot134 bot135 {r}
Lbot_134_135 bot134 bot135 {l}
Rtop_134_164 top134 top164 {r}
Ltop_134_164 top134 top164 {l}
Rbot_134_164 bot134 bot164 {r}
Lbot_134_164 bot134 bot164 {l}
C134 top134 bot134 {c}
Rtop_135_136 top135 top136 {r}
Ltop_135_136 top135 top136 {l}
Rbot_135_136 bot135 bot136 {r}
Lbot_135_136 bot135 bot136 {l}
Rtop_135_165 top135 top165 {r}
Ltop_135_165 top135 top165 {l}
Rbot_135_165 bot135 bot165 {r}
Lbot_135_165 bot135 bot165 {l}
C135 top135 bot135 {c}
Rtop_136_137 top136 top137 {r}
Ltop_136_137 top136 top137 {l}
Rbot_136_137 bot136 bot137 {r}
Lbot_136_137 bot136 bot137 {l}
Rtop_136_166 top136 top166 {r}
Ltop_136_166 top136 top166 {l}
Rbot_136_166 bot136 bot166 {r}
Lbot_136_166 bot136 bot166 {l}
C136 top136 bot136 {c}
Rtop_137_138 top137 top138 {r}
Ltop_137_138 top137 top138 {l}
Rbot_137_138 bot137 bot138 {r}
Lbot_137_138 bot137 bot138 {l}
Rtop_137_167 top137 top167 {r}
Ltop_137_167 top137 top167 {l}
Rbot_137_167 bot137 bot167 {r}
Lbot_137_167 bot137 bot167 {l}
C137 top137 bot137 {c}
Rtop_138_139 top138 top139 {r}
Ltop_138_139 top138 top139 {l}
Rbot_138_139 bot138 bot139 {r}
Lbot_138_139 bot138 bot139 {l}
Rtop_138_168 top138 top168 {r}
Ltop_138_168 top138 top168 {l}
Rbot_138_168 bot138 bot168 {r}
Lbot_138_168 bot138 bot168 {l}
C138 top138 bot138 {c}
Rtop_139_140 top139 top140 {r}
Ltop_139_140 top139 top140 {l}
Rbot_139_140 bot139 bot140 {r}
Lbot_139_140 bot139 bot140 {l}
Rtop_139_169 top139 top169 {r}
Ltop_139_169 top139 top169 {l}
Rbot_139_169 bot139 bot169 {r}
Lbot_139_169 bot139 bot169 {l}
C139 top139 bot139 {c}
Rtop_140_141 top140 top141 {r}
Ltop_140_141 top140 top141 {l}
Rbot_140_141 bot140 bot141 {r}
Lbot_140_141 bot140 bot141 {l}
Rtop_140_170 top140 top170 {r}
Ltop_140_170 top140 top170 {l}
Rbot_140_170 bot140 bot170 {r}
Lbot_140_170 bot140 bot170 {l}
C140 top140 bot140 {c}
Rtop_141_142 top141 top142 {r}
Ltop_141_142 top141 top142 {l}
Rbot_141_142 bot141 bot142 {r}
Lbot_141_142 bot141 bot142 {l}
Rtop_141_171 top141 top171 {r}
Ltop_141_171 top141 top171 {l}
Rbot_141_171 bot141 bot171 {r}
Lbot_141_171 bot141 bot171 {l}
C141 top141 bot141 {c}
Rtop_142_143 top142 top143 {r}
Ltop_142_143 top142 top143 {l}
Rbot_142_143 bot142 bot143 {r}
Lbot_142_143 bot142 bot143 {l}
Rtop_142_172 top142 top172 {r}
Ltop_142_172 top142 top172 {l}
Rbot_142_172 bot142 bot172 {r}
Lbot_142_172 bot142 bot172 {l}
C142 top142 bot142 {c}
Rtop_143_144 top143 top144 {r}
Ltop_143_144 top143 top144 {l}
Rbot_143_144 bot143 bot144 {r}
Lbot_143_144 bot143 bot144 {l}
Rtop_143_173 top143 top173 {r}
Ltop_143_173 top143 top173 {l}
Rbot_143_173 bot143 bot173 {r}
Lbot_143_173 bot143 bot173 {l}
C143 top143 bot143 {c}
Rtop_144_145 top144 top145 {r}
Ltop_144_145 top144 top145 {l}
Rbot_144_145 bot144 bot145 {r}
Lbot_144_145 bot144 bot145 {l}
Rtop_144_174 top144 top174 {r}
Ltop_144_174 top144 top174 {l}
Rbot_144_174 bot144 bot174 {r}
Lbot_144_174 bot144 bot174 {l}
C144 top144 bot144 {c}
Rtop_145_146 top145 top146 {r}
Ltop_145_146 top145 top146 {l}
Rbot_145_146 bot145 bot146 {r}
Lbot_145_146 bot145 bot146 {l}
Rtop_145_175 top145 top175 {r}
Ltop_145_175 top145 top175 {l}
Rbot_145_175 bot145 bot175 {r}
Lbot_145_175 bot145 bot175 {l}
C145 top145 bot145 {c}
Rtop_146_147 top146 top147 {r}
Ltop_146_147 top146 top147 {l}
Rbot_146_147 bot146 bot147 {r}
Lbot_146_147 bot146 bot147 {l}
Rtop_146_176 top146 top176 {r}
Ltop_146_176 top146 top176 {l}
Rbot_146_176 bot146 bot176 {r}
Lbot_146_176 bot146 bot176 {l}
C146 top146 bot146 {c}
Rtop_147_148 top147 top148 {r}
Ltop_147_148 top147 top148 {l}
Rbot_147_148 bot147 bot148 {r}
Lbot_147_148 bot147 bot148 {l}
Rtop_147_177 top147 top177 {r}
Ltop_147_177 top147 top177 {l}
Rbot_147_177 bot147 bot177 {r}
Lbot_147_177 bot147 bot177 {l}
C147 top147 bot147 {c}
Rtop_148_149 top148 top149 {r}
Ltop_148_149 top148 top149 {l}
Rbot_148_149 bot148 bot149 {r}
Lbot_148_149 bot148 bot149 {l}
Rtop_148_178 top148 top178 {r}
Ltop_148_178 top148 top178 {l}
Rbot_148_178 bot148 bot178 {r}
Lbot_148_178 bot148 bot178 {l}
C148 top148 bot148 {c}
Rtop_149_150 top149 top150 {r}
Ltop_149_150 top149 top150 {l}
Rbot_149_150 bot149 bot150 {r}
Lbot_149_150 bot149 bot150 {l}
Rtop_149_179 top149 top179 {r}
Ltop_149_179 top149 top179 {l}
Rbot_149_179 bot149 bot179 {r}
Lbot_149_179 bot149 bot179 {l}
C149 top149 bot149 {c}
Rtop_150_180 top150 top180 {r}
Ltop_150_180 top150 top180 {l}
Rbot_150_180 bot150 bot180 {r}
Lbot_150_180 bot150 bot180 {l}
C150 top150 bot150 {c}
Rtop_151_152 top151 top152 {r}
Ltop_151_152 top151 top152 {l}
Rbot_151_152 bot151 bot152 {r}
Lbot_151_152 bot151 bot152 {l}
Rtop_151_181 top151 top181 {r}
Ltop_151_181 top151 top181 {l}
Rbot_151_181 bot151 bot181 {r}
Lbot_151_181 bot151 bot181 {l}
C151 top151 bot151 {c}
Rtop_152_153 top152 top153 {r}
Ltop_152_153 top152 top153 {l}
Rbot_152_153 bot152 bot153 {r}
Lbot_152_153 bot152 bot153 {l}
Rtop_152_182 top152 top182 {r}
Ltop_152_182 top152 top182 {l}
Rbot_152_182 bot152 bot182 {r}
Lbot_152_182 bot152 bot182 {l}
C152 top152 bot152 {c}
Rtop_153_154 top153 top154 {r}
Ltop_153_154 top153 top154 {l}
Rbot_153_154 bot153 bot154 {r}
Lbot_153_154 bot153 bot154 {l}
Rtop_153_183 top153 top183 {r}
Ltop_153_183 top153 top183 {l}
Rbot_153_183 bot153 bot183 {r}
Lbot_153_183 bot153 bot183 {l}
C153 top153 bot153 {c}
Rtop_154_155 top154 top155 {r}
Ltop_154_155 top154 top155 {l}
Rbot_154_155 bot154 bot155 {r}
Lbot_154_155 bot154 bot155 {l}
Rtop_154_184 top154 top184 {r}
Ltop_154_184 top154 top184 {l}
Rbot_154_184 bot154 bot184 {r}
Lbot_154_184 bot154 bot184 {l}
C154 top154 bot154 {c}
Rtop_155_156 top155 top156 {r}
Ltop_155_156 top155 top156 {l}
Rbot_155_156 bot155 bot156 {r}
Lbot_155_156 bot155 bot156 {l}
Rtop_155_185 top155 top185 {r}
Ltop_155_185 top155 top185 {l}
Rbot_155_185 bot155 bot185 {r}
Lbot_155_185 bot155 bot185 {l}
C155 top155 bot155 {c}
Rtop_156_157 top156 top157 {r}
Ltop_156_157 top156 top157 {l}
Rbot_156_157 bot156 bot157 {r}
Lbot_156_157 bot156 bot157 {l}
Rtop_156_186 top156 top186 {r}
Ltop_156_186 top156 top186 {l}
Rbot_156_186 bot156 bot186 {r}
Lbot_156_186 bot156 bot186 {l}
C156 top156 bot156 {c}
Rtop_157_158 top157 top158 {r}
Ltop_157_158 top157 top158 {l}
Rbot_157_158 bot157 bot158 {r}
Lbot_157_158 bot157 bot158 {l}
Rtop_157_187 top157 top187 {r}
Ltop_157_187 top157 top187 {l}
Rbot_157_187 bot157 bot187 {r}
Lbot_157_187 bot157 bot187 {l}
C157 top157 bot157 {c}
Rtop_158_159 top158 top159 {r}
Ltop_158_159 top158 top159 {l}
Rbot_158_159 bot158 bot159 {r}
Lbot_158_159 bot158 bot159 {l}
Rtop_158_188 top158 top188 {r}
Ltop_158_188 top158 top188 {l}
Rbot_158_188 bot158 bot188 {r}
Lbot_158_188 bot158 bot188 {l}
C158 top158 bot158 {c}
Rtop_159_160 top159 top160 {r}
Ltop_159_160 top159 top160 {l}
Rbot_159_160 bot159 bot160 {r}
Lbot_159_160 bot159 bot160 {l}
Rtop_159_189 top159 top189 {r}
Ltop_159_189 top159 top189 {l}
Rbot_159_189 bot159 bot189 {r}
Lbot_159_189 bot159 bot189 {l}
C159 top159 bot159 {c}
Rtop_160_161 top160 top161 {r}
Ltop_160_161 top160 top161 {l}
Rbot_160_161 bot160 bot161 {r}
Lbot_160_161 bot160 bot161 {l}
Rtop_160_190 top160 top190 {r}
Ltop_160_190 top160 top190 {l}
Rbot_160_190 bot160 bot190 {r}
Lbot_160_190 bot160 bot190 {l}
C160 top160 bot160 {c}
Rtop_161_162 top161 top162 {r}
Ltop_161_162 top161 top162 {l}
Rbot_161_162 bot161 bot162 {r}
Lbot_161_162 bot161 bot162 {l}
Rtop_161_191 top161 top191 {r}
Ltop_161_191 top161 top191 {l}
Rbot_161_191 bot161 bot191 {r}
Lbot_161_191 bot161 bot191 {l}
C161 top161 bot161 {c}
Rtop_162_163 top162 top163 {r}
Ltop_162_163 top162 top163 {l}
Rbot_162_163 bot162 bot163 {r}
Lbot_162_163 bot162 bot163 {l}
Rtop_162_192 top162 top192 {r}
Ltop_162_192 top162 top192 {l}
Rbot_162_192 bot162 bot192 {r}
Lbot_162_192 bot162 bot192 {l}
C162 top162 bot162 {c}
Rtop_163_164 top163 top164 {r}
Ltop_163_164 top163 top164 {l}
Rbot_163_164 bot163 bot164 {r}
Lbot_163_164 bot163 bot164 {l}
Rtop_163_193 top163 top193 {r}
Ltop_163_193 top163 top193 {l}
Rbot_163_193 bot163 bot193 {r}
Lbot_163_193 bot163 bot193 {l}
C163 top163 bot163 {c}
Rtop_164_165 top164 top165 {r}
Ltop_164_165 top164 top165 {l}
Rbot_164_165 bot164 bot165 {r}
Lbot_164_165 bot164 bot165 {l}
Rtop_164_194 top164 top194 {r}
Ltop_164_194 top164 top194 {l}
Rbot_164_194 bot164 bot194 {r}
Lbot_164_194 bot164 bot194 {l}
C164 top164 bot164 {c}
Rtop_165_166 top165 top166 {r}
Ltop_165_166 top165 top166 {l}
Rbot_165_166 bot165 bot166 {r}
Lbot_165_166 bot165 bot166 {l}
Rtop_165_195 top165 top195 {r}
Ltop_165_195 top165 top195 {l}
Rbot_165_195 bot165 bot195 {r}
Lbot_165_195 bot165 bot195 {l}
C165 top165 bot165 {c}
Rtop_166_167 top166 top167 {r}
Ltop_166_167 top166 top167 {l}
Rbot_166_167 bot166 bot167 {r}
Lbot_166_167 bot166 bot167 {l}
Rtop_166_196 top166 top196 {r}
Ltop_166_196 top166 top196 {l}
Rbot_166_196 bot166 bot196 {r}
Lbot_166_196 bot166 bot196 {l}
C166 top166 bot166 {c}
Rtop_167_168 top167 top168 {r}
Ltop_167_168 top167 top168 {l}
Rbot_167_168 bot167 bot168 {r}
Lbot_167_168 bot167 bot168 {l}
Rtop_167_197 top167 top197 {r}
Ltop_167_197 top167 top197 {l}
Rbot_167_197 bot167 bot197 {r}
Lbot_167_197 bot167 bot197 {l}
C167 top167 bot167 {c}
Rtop_168_169 top168 top169 {r}
Ltop_168_169 top168 top169 {l}
Rbot_168_169 bot168 bot169 {r}
Lbot_168_169 bot168 bot169 {l}
Rtop_168_198 top168 top198 {r}
Ltop_168_198 top168 top198 {l}
Rbot_168_198 bot168 bot198 {r}
Lbot_168_198 bot168 bot198 {l}
C168 top168 bot168 {c}
Rtop_169_170 top169 top170 {r}
Ltop_169_170 top169 top170 {l}
Rbot_169_170 bot169 bot170 {r}
Lbot_169_170 bot169 bot170 {l}
Rtop_169_199 top169 top199 {r}
Ltop_169_199 top169 top199 {l}
Rbot_169_199 bot169 bot199 {r}
Lbot_169_199 bot169 bot199 {l}
C169 top169 bot169 {c}
Rtop_170_171 top170 top171 {r}
Ltop_170_171 top170 top171 {l}
Rbot_170_171 bot170 bot171 {r}
Lbot_170_171 bot170 bot171 {l}
Rtop_170_200 top170 top200 {r}
Ltop_170_200 top170 top200 {l}
Rbot_170_200 bot170 bot200 {r}
Lbot_170_200 bot170 bot200 {l}
C170 top170 bot170 {c}
Rtop_171_172 top171 top172 {r}
Ltop_171_172 top171 top172 {l}
Rbot_171_172 bot171 bot172 {r}
Lbot_171_172 bot171 bot172 {l}
Rtop_171_201 top171 top201 {r}
Ltop_171_201 top171 top201 {l}
Rbot_171_201 bot171 bot201 {r}
Lbot_171_201 bot171 bot201 {l}
C171 top171 bot171 {c}
Rtop_172_173 top172 top173 {r}
Ltop_172_173 top172 top173 {l}
Rbot_172_173 bot172 bot173 {r}
Lbot_172_173 bot172 bot173 {l}
Rtop_172_202 top172 top202 {r}
Ltop_172_202 top172 top202 {l}
Rbot_172_202 bot172 bot202 {r}
Lbot_172_202 bot172 bot202 {l}
C172 top172 bot172 {c}
Rtop_173_174 top173 top174 {r}
Ltop_173_174 top173 top174 {l}
Rbot_173_174 bot173 bot174 {r}
Lbot_173_174 bot173 bot174 {l}
Rtop_173_203 top173 top203 {r}
Ltop_173_203 top173 top203 {l}
Rbot_173_203 bot173 bot203 {r}
Lbot_173_203 bot173 bot203 {l}
C173 top173 bot173 {c}
Rtop_174_175 top174 top175 {r}
Ltop_174_175 top174 top175 {l}
Rbot_174_175 bot174 bot175 {r}
Lbot_174_175 bot174 bot175 {l}
Rtop_174_204 top174 top204 {r}
Ltop_174_204 top174 top204 {l}
Rbot_174_204 bot174 bot204 {r}
Lbot_174_204 bot174 bot204 {l}
C174 top174 bot174 {c}
Rtop_175_176 top175 top176 {r}
Ltop_175_176 top175 top176 {l}
Rbot_175_176 bot175 bot176 {r}
Lbot_175_176 bot175 bot176 {l}
Rtop_175_205 top175 top205 {r}
Ltop_175_205 top175 top205 {l}
Rbot_175_205 bot175 bot205 {r}
Lbot_175_205 bot175 bot205 {l}
C175 top175 bot175 {c}
Rtop_176_177 top176 top177 {r}
Ltop_176_177 top176 top177 {l}
Rbot_176_177 bot176 bot177 {r}
Lbot_176_177 bot176 bot177 {l}
Rtop_176_206 top176 top206 {r}
Ltop_176_206 top176 top206 {l}
Rbot_176_206 bot176 bot206 {r}
Lbot_176_206 bot176 bot206 {l}
C176 top176 bot176 {c}
Rtop_177_178 top177 top178 {r}
Ltop_177_178 top177 top178 {l}
Rbot_177_178 bot177 bot178 {r}
Lbot_177_178 bot177 bot178 {l}
Rtop_177_207 top177 top207 {r}
Ltop_177_207 top177 top207 {l}
Rbot_177_207 bot177 bot207 {r}
Lbot_177_207 bot177 bot207 {l}
C177 top177 bot177 {c}
Rtop_178_179 top178 top179 {r}
Ltop_178_179 top178 top179 {l}
Rbot_178_179 bot178 bot179 {r}
Lbot_178_179 bot178 bot179 {l}
Rtop_178_208 top178 top208 {r}
Ltop_178_208 top178 top208 {l}
Rbot_178_208 bot178 bot208 {r}
Lbot_178_208 bot178 bot208 {l}
C178 top178 bot178 {c}
Rtop_179_180 top179 top180 {r}
Ltop_179_180 top179 top180 {l}
Rbot_179_180 bot179 bot180 {r}
Lbot_179_180 bot179 bot180 {l}
Rtop_179_209 top179 top209 {r}
Ltop_179_209 top179 top209 {l}
Rbot_179_209 bot179 bot209 {r}
Lbot_179_209 bot179 bot209 {l}
C179 top179 bot179 {c}
Rtop_180_210 top180 top210 {r}
Ltop_180_210 top180 top210 {l}
Rbot_180_210 bot180 bot210 {r}
Lbot_180_210 bot180 bot210 {l}
C180 top180 bot180 {c}
Rtop_181_182 top181 top182 {r}
Ltop_181_182 top181 top182 {l}
Rbot_181_182 bot181 bot182 {r}
Lbot_181_182 bot181 bot182 {l}
Rtop_181_211 top181 top211 {r}
Ltop_181_211 top181 top211 {l}
Rbot_181_211 bot181 bot211 {r}
Lbot_181_211 bot181 bot211 {l}
C181 top181 bot181 {c}
Rtop_182_183 top182 top183 {r}
Ltop_182_183 top182 top183 {l}
Rbot_182_183 bot182 bot183 {r}
Lbot_182_183 bot182 bot183 {l}
Rtop_182_212 top182 top212 {r}
Ltop_182_212 top182 top212 {l}
Rbot_182_212 bot182 bot212 {r}
Lbot_182_212 bot182 bot212 {l}
C182 top182 bot182 {c}
Rtop_183_184 top183 top184 {r}
Ltop_183_184 top183 top184 {l}
Rbot_183_184 bot183 bot184 {r}
Lbot_183_184 bot183 bot184 {l}
Rtop_183_213 top183 top213 {r}
Ltop_183_213 top183 top213 {l}
Rbot_183_213 bot183 bot213 {r}
Lbot_183_213 bot183 bot213 {l}
C183 top183 bot183 {c}
Rtop_184_185 top184 top185 {r}
Ltop_184_185 top184 top185 {l}
Rbot_184_185 bot184 bot185 {r}
Lbot_184_185 bot184 bot185 {l}
Rtop_184_214 top184 top214 {r}
Ltop_184_214 top184 top214 {l}
Rbot_184_214 bot184 bot214 {r}
Lbot_184_214 bot184 bot214 {l}
C184 top184 bot184 {c}
Rtop_185_186 top185 top186 {r}
Ltop_185_186 top185 top186 {l}
Rbot_185_186 bot185 bot186 {r}
Lbot_185_186 bot185 bot186 {l}
Rtop_185_215 top185 top215 {r}
Ltop_185_215 top185 top215 {l}
Rbot_185_215 bot185 bot215 {r}
Lbot_185_215 bot185 bot215 {l}
C185 top185 bot185 {c}
Rtop_186_187 top186 top187 {r}
Ltop_186_187 top186 top187 {l}
Rbot_186_187 bot186 bot187 {r}
Lbot_186_187 bot186 bot187 {l}
Rtop_186_216 top186 top216 {r}
Ltop_186_216 top186 top216 {l}
Rbot_186_216 bot186 bot216 {r}
Lbot_186_216 bot186 bot216 {l}
C186 top186 bot186 {c}
Rtop_187_188 top187 top188 {r}
Ltop_187_188 top187 top188 {l}
Rbot_187_188 bot187 bot188 {r}
Lbot_187_188 bot187 bot188 {l}
Rtop_187_217 top187 top217 {r}
Ltop_187_217 top187 top217 {l}
Rbot_187_217 bot187 bot217 {r}
Lbot_187_217 bot187 bot217 {l}
C187 top187 bot187 {c}
Rtop_188_189 top188 top189 {r}
Ltop_188_189 top188 top189 {l}
Rbot_188_189 bot188 bot189 {r}
Lbot_188_189 bot188 bot189 {l}
Rtop_188_218 top188 top218 {r}
Ltop_188_218 top188 top218 {l}
Rbot_188_218 bot188 bot218 {r}
Lbot_188_218 bot188 bot218 {l}
C188 top188 bot188 {c}
Rtop_189_190 top189 top190 {r}
Ltop_189_190 top189 top190 {l}
Rbot_189_190 bot189 bot190 {r}
Lbot_189_190 bot189 bot190 {l}
Rtop_189_219 top189 top219 {r}
Ltop_189_219 top189 top219 {l}
Rbot_189_219 bot189 bot219 {r}
Lbot_189_219 bot189 bot219 {l}
C189 top189 bot189 {c}
Rtop_190_191 top190 top191 {r}
Ltop_190_191 top190 top191 {l}
Rbot_190_191 bot190 bot191 {r}
Lbot_190_191 bot190 bot191 {l}
Rtop_190_220 top190 top220 {r}
Ltop_190_220 top190 top220 {l}
Rbot_190_220 bot190 bot220 {r}
Lbot_190_220 bot190 bot220 {l}
C190 top190 bot190 {c}
Rtop_191_192 top191 top192 {r}
Ltop_191_192 top191 top192 {l}
Rbot_191_192 bot191 bot192 {r}
Lbot_191_192 bot191 bot192 {l}
Rtop_191_221 top191 top221 {r}
Ltop_191_221 top191 top221 {l}
Rbot_191_221 bot191 bot221 {r}
Lbot_191_221 bot191 bot221 {l}
C191 top191 bot191 {c}
Rtop_192_193 top192 top193 {r}
Ltop_192_193 top192 top193 {l}
Rbot_192_193 bot192 bot193 {r}
Lbot_192_193 bot192 bot193 {l}
Rtop_192_222 top192 top222 {r}
Ltop_192_222 top192 top222 {l}
Rbot_192_222 bot192 bot222 {r}
Lbot_192_222 bot192 bot222 {l}
C192 top192 bot192 {c}
Rtop_193_194 top193 top194 {r}
Ltop_193_194 top193 top194 {l}
Rbot_193_194 bot193 bot194 {r}
Lbot_193_194 bot193 bot194 {l}
Rtop_193_223 top193 top223 {r}
Ltop_193_223 top193 top223 {l}
Rbot_193_223 bot193 bot223 {r}
Lbot_193_223 bot193 bot223 {l}
C193 top193 bot193 {c}
Rtop_194_195 top194 top195 {r}
Ltop_194_195 top194 top195 {l}
Rbot_194_195 bot194 bot195 {r}
Lbot_194_195 bot194 bot195 {l}
Rtop_194_224 top194 top224 {r}
Ltop_194_224 top194 top224 {l}
Rbot_194_224 bot194 bot224 {r}
Lbot_194_224 bot194 bot224 {l}
C194 top194 bot194 {c}
Rtop_195_196 top195 top196 {r}
Ltop_195_196 top195 top196 {l}
Rbot_195_196 bot195 bot196 {r}
Lbot_195_196 bot195 bot196 {l}
Rtop_195_225 top195 top225 {r}
Ltop_195_225 top195 top225 {l}
Rbot_195_225 bot195 bot225 {r}
Lbot_195_225 bot195 bot225 {l}
C195 top195 bot195 {c}
Rtop_196_197 top196 top197 {r}
Ltop_196_197 top196 top197 {l}
Rbot_196_197 bot196 bot197 {r}
Lbot_196_197 bot196 bot197 {l}
Rtop_196_226 top196 top226 {r}
Ltop_196_226 top196 top226 {l}
Rbot_196_226 bot196 bot226 {r}
Lbot_196_226 bot196 bot226 {l}
C196 top196 bot196 {c}
Rtop_197_198 top197 top198 {r}
Ltop_197_198 top197 top198 {l}
Rbot_197_198 bot197 bot198 {r}
Lbot_197_198 bot197 bot198 {l}
Rtop_197_227 top197 top227 {r}
Ltop_197_227 top197 top227 {l}
Rbot_197_227 bot197 bot227 {r}
Lbot_197_227 bot197 bot227 {l}
C197 top197 bot197 {c}
Rtop_198_199 top198 top199 {r}
Ltop_198_199 top198 top199 {l}
Rbot_198_199 bot198 bot199 {r}
Lbot_198_199 bot198 bot199 {l}
Rtop_198_228 top198 top228 {r}
Ltop_198_228 top198 top228 {l}
Rbot_198_228 bot198 bot228 {r}
Lbot_198_228 bot198 bot228 {l}
C198 top198 bot198 {c}
Rtop_199_200 top199 top200 {r}
Ltop_199_200 top199 top200 {l}
Rbot_199_200 bot199 bot200 {r}
Lbot_199_200 bot199 bot200 {l}
Rtop_199_229 top199 top229 {r}
Ltop_199_229 top199 top229 {l}
Rbot_199_229 bot199 bot229 {r}
Lbot_199_229 bot199 bot229 {l}
C199 top199 bot199 {c}
Rtop_200_201 top200 top201 {r}
Ltop_200_201 top200 top201 {l}
Rbot_200_201 bot200 bot201 {r}
Lbot_200_201 bot200 bot201 {l}
Rtop_200_230 top200 top230 {r}
Ltop_200_230 top200 top230 {l}
Rbot_200_230 bot200 bot230 {r}
Lbot_200_230 bot200 bot230 {l}
C200 top200 bot200 {c}
Rtop_201_202 top201 top202 {r}
Ltop_201_202 top201 top202 {l}
Rbot_201_202 bot201 bot202 {r}
Lbot_201_202 bot201 bot202 {l}
Rtop_201_231 top201 top231 {r}
Ltop_201_231 top201 top231 {l}
Rbot_201_231 bot201 bot231 {r}
Lbot_201_231 bot201 bot231 {l}
C201 top201 bot201 {c}
Rtop_202_203 top202 top203 {r}
Ltop_202_203 top202 top203 {l}
Rbot_202_203 bot202 bot203 {r}
Lbot_202_203 bot202 bot203 {l}
Rtop_202_232 top202 top232 {r}
Ltop_202_232 top202 top232 {l}
Rbot_202_232 bot202 bot232 {r}
Lbot_202_232 bot202 bot232 {l}
C202 top202 bot202 {c}
Rtop_203_204 top203 top204 {r}
Ltop_203_204 top203 top204 {l}
Rbot_203_204 bot203 bot204 {r}
Lbot_203_204 bot203 bot204 {l}
Rtop_203_233 top203 top233 {r}
Ltop_203_233 top203 top233 {l}
Rbot_203_233 bot203 bot233 {r}
Lbot_203_233 bot203 bot233 {l}
C203 top203 bot203 {c}
Rtop_204_205 top204 top205 {r}
Ltop_204_205 top204 top205 {l}
Rbot_204_205 bot204 bot205 {r}
Lbot_204_205 bot204 bot205 {l}
Rtop_204_234 top204 top234 {r}
Ltop_204_234 top204 top234 {l}
Rbot_204_234 bot204 bot234 {r}
Lbot_204_234 bot204 bot234 {l}
C204 top204 bot204 {c}
Rtop_205_206 top205 top206 {r}
Ltop_205_206 top205 top206 {l}
Rbot_205_206 bot205 bot206 {r}
Lbot_205_206 bot205 bot206 {l}
Rtop_205_235 top205 top235 {r}
Ltop_205_235 top205 top235 {l}
Rbot_205_235 bot205 bot235 {r}
Lbot_205_235 bot205 bot235 {l}
C205 top205 bot205 {c}
Rtop_206_207 top206 top207 {r}
Ltop_206_207 top206 top207 {l}
Rbot_206_207 bot206 bot207 {r}
Lbot_206_207 bot206 bot207 {l}
Rtop_206_236 top206 top236 {r}
Ltop_206_236 top206 top236 {l}
Rbot_206_236 bot206 bot236 {r}
Lbot_206_236 bot206 bot236 {l}
C206 top206 bot206 {c}
Rtop_207_208 top207 top208 {r}
Ltop_207_208 top207 top208 {l}
Rbot_207_208 bot207 bot208 {r}
Lbot_207_208 bot207 bot208 {l}
Rtop_207_237 top207 top237 {r}
Ltop_207_237 top207 top237 {l}
Rbot_207_237 bot207 bot237 {r}
Lbot_207_237 bot207 bot237 {l}
C207 top207 bot207 {c}
Rtop_208_209 top208 top209 {r}
Ltop_208_209 top208 top209 {l}
Rbot_208_209 bot208 bot209 {r}
Lbot_208_209 bot208 bot209 {l}
Rtop_208_238 top208 top238 {r}
Ltop_208_238 top208 top238 {l}
Rbot_208_238 bot208 bot238 {r}
Lbot_208_238 bot208 bot238 {l}
C208 top208 bot208 {c}
Rtop_209_210 top209 top210 {r}
Ltop_209_210 top209 top210 {l}
Rbot_209_210 bot209 bot210 {r}
Lbot_209_210 bot209 bot210 {l}
Rtop_209_239 top209 top239 {r}
Ltop_209_239 top209 top239 {l}
Rbot_209_239 bot209 bot239 {r}
Lbot_209_239 bot209 bot239 {l}
C209 top209 bot209 {c}
Rtop_210_240 top210 top240 {r}
Ltop_210_240 top210 top240 {l}
Rbot_210_240 bot210 bot240 {r}
Lbot_210_240 bot210 bot240 {l}
C210 top210 bot210 {c}
Rtop_211_212 top211 top212 {r}
Ltop_211_212 top211 top212 {l}
Rbot_211_212 bot211 bot212 {r}
Lbot_211_212 bot211 bot212 {l}
Rtop_211_241 top211 top241 {r}
Ltop_211_241 top211 top241 {l}
Rbot_211_241 bot211 bot241 {r}
Lbot_211_241 bot211 bot241 {l}
C211 top211 bot211 {c}
Rtop_212_213 top212 top213 {r}
Ltop_212_213 top212 top213 {l}
Rbot_212_213 bot212 bot213 {r}
Lbot_212_213 bot212 bot213 {l}
Rtop_212_242 top212 top242 {r}
Ltop_212_242 top212 top242 {l}
Rbot_212_242 bot212 bot242 {r}
Lbot_212_242 bot212 bot242 {l}
C212 top212 bot212 {c}
Rtop_213_214 top213 top214 {r}
Ltop_213_214 top213 top214 {l}
Rbot_213_214 bot213 bot214 {r}
Lbot_213_214 bot213 bot214 {l}
Rtop_213_243 top213 top243 {r}
Ltop_213_243 top213 top243 {l}
Rbot_213_243 bot213 bot243 {r}
Lbot_213_243 bot213 bot243 {l}
C213 top213 bot213 {c}
Rtop_214_215 top214 top215 {r}
Ltop_214_215 top214 top215 {l}
Rbot_214_215 bot214 bot215 {r}
Lbot_214_215 bot214 bot215 {l}
Rtop_214_244 top214 top244 {r}
Ltop_214_244 top214 top244 {l}
Rbot_214_244 bot214 bot244 {r}
Lbot_214_244 bot214 bot244 {l}
C214 top214 bot214 {c}
Rtop_215_216 top215 top216 {r}
Ltop_215_216 top215 top216 {l}
Rbot_215_216 bot215 bot216 {r}
Lbot_215_216 bot215 bot216 {l}
Rtop_215_245 top215 top245 {r}
Ltop_215_245 top215 top245 {l}
Rbot_215_245 bot215 bot245 {r}
Lbot_215_245 bot215 bot245 {l}
C215 top215 bot215 {c}
Rtop_216_217 top216 top217 {r}
Ltop_216_217 top216 top217 {l}
Rbot_216_217 bot216 bot217 {r}
Lbot_216_217 bot216 bot217 {l}
Rtop_216_246 top216 top246 {r}
Ltop_216_246 top216 top246 {l}
Rbot_216_246 bot216 bot246 {r}
Lbot_216_246 bot216 bot246 {l}
C216 top216 bot216 {c}
Rtop_217_218 top217 top218 {r}
Ltop_217_218 top217 top218 {l}
Rbot_217_218 bot217 bot218 {r}
Lbot_217_218 bot217 bot218 {l}
Rtop_217_247 top217 top247 {r}
Ltop_217_247 top217 top247 {l}
Rbot_217_247 bot217 bot247 {r}
Lbot_217_247 bot217 bot247 {l}
C217 top217 bot217 {c}
Rtop_218_219 top218 top219 {r}
Ltop_218_219 top218 top219 {l}
Rbot_218_219 bot218 bot219 {r}
Lbot_218_219 bot218 bot219 {l}
Rtop_218_248 top218 top248 {r}
Ltop_218_248 top218 top248 {l}
Rbot_218_248 bot218 bot248 {r}
Lbot_218_248 bot218 bot248 {l}
C218 top218 bot218 {c}
Rtop_219_220 top219 top220 {r}
Ltop_219_220 top219 top220 {l}
Rbot_219_220 bot219 bot220 {r}
Lbot_219_220 bot219 bot220 {l}
Rtop_219_249 top219 top249 {r}
Ltop_219_249 top219 top249 {l}
Rbot_219_249 bot219 bot249 {r}
Lbot_219_249 bot219 bot249 {l}
C219 top219 bot219 {c}
Rtop_220_221 top220 top221 {r}
Ltop_220_221 top220 top221 {l}
Rbot_220_221 bot220 bot221 {r}
Lbot_220_221 bot220 bot221 {l}
Rtop_220_250 top220 top250 {r}
Ltop_220_250 top220 top250 {l}
Rbot_220_250 bot220 bot250 {r}
Lbot_220_250 bot220 bot250 {l}
C220 top220 bot220 {c}
Rtop_221_222 top221 top222 {r}
Ltop_221_222 top221 top222 {l}
Rbot_221_222 bot221 bot222 {r}
Lbot_221_222 bot221 bot222 {l}
Rtop_221_251 top221 top251 {r}
Ltop_221_251 top221 top251 {l}
Rbot_221_251 bot221 bot251 {r}
Lbot_221_251 bot221 bot251 {l}
C221 top221 bot221 {c}
Rtop_222_223 top222 top223 {r}
Ltop_222_223 top222 top223 {l}
Rbot_222_223 bot222 bot223 {r}
Lbot_222_223 bot222 bot223 {l}
Rtop_222_252 top222 top252 {r}
Ltop_222_252 top222 top252 {l}
Rbot_222_252 bot222 bot252 {r}
Lbot_222_252 bot222 bot252 {l}
C222 top222 bot222 {c}
Rtop_223_224 top223 top224 {r}
Ltop_223_224 top223 top224 {l}
Rbot_223_224 bot223 bot224 {r}
Lbot_223_224 bot223 bot224 {l}
Rtop_223_253 top223 top253 {r}
Ltop_223_253 top223 top253 {l}
Rbot_223_253 bot223 bot253 {r}
Lbot_223_253 bot223 bot253 {l}
C223 top223 bot223 {c}
Rtop_224_225 top224 top225 {r}
Ltop_224_225 top224 top225 {l}
Rbot_224_225 bot224 bot225 {r}
Lbot_224_225 bot224 bot225 {l}
Rtop_224_254 top224 top254 {r}
Ltop_224_254 top224 top254 {l}
Rbot_224_254 bot224 bot254 {r}
Lbot_224_254 bot224 bot254 {l}
C224 top224 bot224 {c}
Rtop_225_226 top225 top226 {r}
Ltop_225_226 top225 top226 {l}
Rbot_225_226 bot225 bot226 {r}
Lbot_225_226 bot225 bot226 {l}
Rtop_225_255 top225 top255 {r}
Ltop_225_255 top225 top255 {l}
Rbot_225_255 bot225 bot255 {r}
Lbot_225_255 bot225 bot255 {l}
C225 top225 bot225 {c}
Rtop_226_227 top226 top227 {r}
Ltop_226_227 top226 top227 {l}
Rbot_226_227 bot226 bot227 {r}
Lbot_226_227 bot226 bot227 {l}
Rtop_226_256 top226 top256 {r}
Ltop_226_256 top226 top256 {l}
Rbot_226_256 bot226 bot256 {r}
Lbot_226_256 bot226 bot256 {l}
C226 top226 bot226 {c}
Rtop_227_228 top227 top228 {r}
Ltop_227_228 top227 top228 {l}
Rbot_227_228 bot227 bot228 {r}
Lbot_227_228 bot227 bot228 {l}
Rtop_227_257 top227 top257 {r}
Ltop_227_257 top227 top257 {l}
Rbot_227_257 bot227 bot257 {r}
Lbot_227_257 bot227 bot257 {l}
C227 top227 bot227 {c}
Rtop_228_229 top228 top229 {r}
Ltop_228_229 top228 top229 {l}
Rbot_228_229 bot228 bot229 {r}
Lbot_228_229 bot228 bot229 {l}
Rtop_228_258 top228 top258 {r}
Ltop_228_258 top228 top258 {l}
Rbot_228_258 bot228 bot258 {r}
Lbot_228_258 bot228 bot258 {l}
C228 top228 bot228 {c}
Rtop_229_230 top229 top230 {r}
Ltop_229_230 top229 top230 {l}
Rbot_229_230 bot229 bot230 {r}
Lbot_229_230 bot229 bot230 {l}
Rtop_229_259 top229 top259 {r}
Ltop_229_259 top229 top259 {l}
Rbot_229_259 bot229 bot259 {r}
Lbot_229_259 bot229 bot259 {l}
C229 top229 bot229 {c}
Rtop_230_231 top230 top231 {r}
Ltop_230_231 top230 top231 {l}
Rbot_230_231 bot230 bot231 {r}
Lbot_230_231 bot230 bot231 {l}
Rtop_230_260 top230 top260 {r}
Ltop_230_260 top230 top260 {l}
Rbot_230_260 bot230 bot260 {r}
Lbot_230_260 bot230 bot260 {l}
C230 top230 bot230 {c}
Rtop_231_232 top231 top232 {r}
Ltop_231_232 top231 top232 {l}
Rbot_231_232 bot231 bot232 {r}
Lbot_231_232 bot231 bot232 {l}
Rtop_231_261 top231 top261 {r}
Ltop_231_261 top231 top261 {l}
Rbot_231_261 bot231 bot261 {r}
Lbot_231_261 bot231 bot261 {l}
C231 top231 bot231 {c}
Rtop_232_233 top232 top233 {r}
Ltop_232_233 top232 top233 {l}
Rbot_232_233 bot232 bot233 {r}
Lbot_232_233 bot232 bot233 {l}
Rtop_232_262 top232 top262 {r}
Ltop_232_262 top232 top262 {l}
Rbot_232_262 bot232 bot262 {r}
Lbot_232_262 bot232 bot262 {l}
C232 top232 bot232 {c}
Rtop_233_234 top233 top234 {r}
Ltop_233_234 top233 top234 {l}
Rbot_233_234 bot233 bot234 {r}
Lbot_233_234 bot233 bot234 {l}
Rtop_233_263 top233 top263 {r}
Ltop_233_263 top233 top263 {l}
Rbot_233_263 bot233 bot263 {r}
Lbot_233_263 bot233 bot263 {l}
C233 top233 bot233 {c}
Rtop_234_235 top234 top235 {r}
Ltop_234_235 top234 top235 {l}
Rbot_234_235 bot234 bot235 {r}
Lbot_234_235 bot234 bot235 {l}
Rtop_234_264 top234 top264 {r}
Ltop_234_264 top234 top264 {l}
Rbot_234_264 bot234 bot264 {r}
Lbot_234_264 bot234 bot264 {l}
C234 top234 bot234 {c}
Rtop_235_236 top235 top236 {r}
Ltop_235_236 top235 top236 {l}
Rbot_235_236 bot235 bot236 {r}
Lbot_235_236 bot235 bot236 {l}
Rtop_235_265 top235 top265 {r}
Ltop_235_265 top235 top265 {l}
Rbot_235_265 bot235 bot265 {r}
Lbot_235_265 bot235 bot265 {l}
C235 top235 bot235 {c}
Rtop_236_237 top236 top237 {r}
Ltop_236_237 top236 top237 {l}
Rbot_236_237 bot236 bot237 {r}
Lbot_236_237 bot236 bot237 {l}
Rtop_236_266 top236 top266 {r}
Ltop_236_266 top236 top266 {l}
Rbot_236_266 bot236 bot266 {r}
Lbot_236_266 bot236 bot266 {l}
C236 top236 bot236 {c}
Rtop_237_238 top237 top238 {r}
Ltop_237_238 top237 top238 {l}
Rbot_237_238 bot237 bot238 {r}
Lbot_237_238 bot237 bot238 {l}
Rtop_237_267 top237 top267 {r}
Ltop_237_267 top237 top267 {l}
Rbot_237_267 bot237 bot267 {r}
Lbot_237_267 bot237 bot267 {l}
C237 top237 bot237 {c}
Rtop_238_239 top238 top239 {r}
Ltop_238_239 top238 top239 {l}
Rbot_238_239 bot238 bot239 {r}
Lbot_238_239 bot238 bot239 {l}
Rtop_238_268 top238 top268 {r}
Ltop_238_268 top238 top268 {l}
Rbot_238_268 bot238 bot268 {r}
Lbot_238_268 bot238 bot268 {l}
C238 top238 bot238 {c}
Rtop_239_240 top239 top240 {r}
Ltop_239_240 top239 top240 {l}
Rbot_239_240 bot239 bot240 {r}
Lbot_239_240 bot239 bot240 {l}
Rtop_239_269 top239 top269 {r}
Ltop_239_269 top239 top269 {l}
Rbot_239_269 bot239 bot269 {r}
Lbot_239_269 bot239 bot269 {l}
C239 top239 bot239 {c}
Rtop_240_270 top240 top270 {r}
Ltop_240_270 top240 top270 {l}
Rbot_240_270 bot240 bot270 {r}
Lbot_240_270 bot240 bot270 {l}
C240 top240 bot240 {c}
Rtop_241_242 top241 top242 {r}
Ltop_241_242 top241 top242 {l}
Rbot_241_242 bot241 bot242 {r}
Lbot_241_242 bot241 bot242 {l}
Rtop_241_271 top241 top271 {r}
Ltop_241_271 top241 top271 {l}
Rbot_241_271 bot241 bot271 {r}
Lbot_241_271 bot241 bot271 {l}
C241 top241 bot241 {c}
Rtop_242_243 top242 top243 {r}
Ltop_242_243 top242 top243 {l}
Rbot_242_243 bot242 bot243 {r}
Lbot_242_243 bot242 bot243 {l}
Rtop_242_272 top242 top272 {r}
Ltop_242_272 top242 top272 {l}
Rbot_242_272 bot242 bot272 {r}
Lbot_242_272 bot242 bot272 {l}
C242 top242 bot242 {c}
Rtop_243_244 top243 top244 {r}
Ltop_243_244 top243 top244 {l}
Rbot_243_244 bot243 bot244 {r}
Lbot_243_244 bot243 bot244 {l}
Rtop_243_273 top243 top273 {r}
Ltop_243_273 top243 top273 {l}
Rbot_243_273 bot243 bot273 {r}
Lbot_243_273 bot243 bot273 {l}
C243 top243 bot243 {c}
Rtop_244_245 top244 top245 {r}
Ltop_244_245 top244 top245 {l}
Rbot_244_245 bot244 bot245 {r}
Lbot_244_245 bot244 bot245 {l}
Rtop_244_274 top244 top274 {r}
Ltop_244_274 top244 top274 {l}
Rbot_244_274 bot244 bot274 {r}
Lbot_244_274 bot244 bot274 {l}
C244 top244 bot244 {c}
Rtop_245_246 top245 top246 {r}
Ltop_245_246 top245 top246 {l}
Rbot_245_246 bot245 bot246 {r}
Lbot_245_246 bot245 bot246 {l}
Rtop_245_275 top245 top275 {r}
Ltop_245_275 top245 top275 {l}
Rbot_245_275 bot245 bot275 {r}
Lbot_245_275 bot245 bot275 {l}
C245 top245 bot245 {c}
Rtop_246_247 top246 top247 {r}
Ltop_246_247 top246 top247 {l}
Rbot_246_247 bot246 bot247 {r}
Lbot_246_247 bot246 bot247 {l}
Rtop_246_276 top246 top276 {r}
Ltop_246_276 top246 top276 {l}
Rbot_246_276 bot246 bot276 {r}
Lbot_246_276 bot246 bot276 {l}
C246 top246 bot246 {c}
Rtop_247_248 top247 top248 {r}
Ltop_247_248 top247 top248 {l}
Rbot_247_248 bot247 bot248 {r}
Lbot_247_248 bot247 bot248 {l}
Rtop_247_277 top247 top277 {r}
Ltop_247_277 top247 top277 {l}
Rbot_247_277 bot247 bot277 {r}
Lbot_247_277 bot247 bot277 {l}
C247 top247 bot247 {c}
Rtop_248_249 top248 top249 {r}
Ltop_248_249 top248 top249 {l}
Rbot_248_249 bot248 bot249 {r}
Lbot_248_249 bot248 bot249 {l}
Rtop_248_278 top248 top278 {r}
Ltop_248_278 top248 top278 {l}
Rbot_248_278 bot248 bot278 {r}
Lbot_248_278 bot248 bot278 {l}
C248 top248 bot248 {c}
Rtop_249_250 top249 top250 {r}
Ltop_249_250 top249 top250 {l}
Rbot_249_250 bot249 bot250 {r}
Lbot_249_250 bot249 bot250 {l}
Rtop_249_279 top249 top279 {r}
Ltop_249_279 top249 top279 {l}
Rbot_249_279 bot249 bot279 {r}
Lbot_249_279 bot249 bot279 {l}
C249 top249 bot249 {c}
Rtop_250_251 top250 top251 {r}
Ltop_250_251 top250 top251 {l}
Rbot_250_251 bot250 bot251 {r}
Lbot_250_251 bot250 bot251 {l}
Rtop_250_280 top250 top280 {r}
Ltop_250_280 top250 top280 {l}
Rbot_250_280 bot250 bot280 {r}
Lbot_250_280 bot250 bot280 {l}
C250 top250 bot250 {c}
Rtop_251_252 top251 top252 {r}
Ltop_251_252 top251 top252 {l}
Rbot_251_252 bot251 bot252 {r}
Lbot_251_252 bot251 bot252 {l}
Rtop_251_281 top251 top281 {r}
Ltop_251_281 top251 top281 {l}
Rbot_251_281 bot251 bot281 {r}
Lbot_251_281 bot251 bot281 {l}
C251 top251 bot251 {c}
Rtop_252_253 top252 top253 {r}
Ltop_252_253 top252 top253 {l}
Rbot_252_253 bot252 bot253 {r}
Lbot_252_253 bot252 bot253 {l}
Rtop_252_282 top252 top282 {r}
Ltop_252_282 top252 top282 {l}
Rbot_252_282 bot252 bot282 {r}
Lbot_252_282 bot252 bot282 {l}
C252 top252 bot252 {c}
Rtop_253_254 top253 top254 {r}
Ltop_253_254 top253 top254 {l}
Rbot_253_254 bot253 bot254 {r}
Lbot_253_254 bot253 bot254 {l}
Rtop_253_283 top253 top283 {r}
Ltop_253_283 top253 top283 {l}
Rbot_253_283 bot253 bot283 {r}
Lbot_253_283 bot253 bot283 {l}
C253 top253 bot253 {c}
Rtop_254_255 top254 top255 {r}
Ltop_254_255 top254 top255 {l}
Rbot_254_255 bot254 bot255 {r}
Lbot_254_255 bot254 bot255 {l}
Rtop_254_284 top254 top284 {r}
Ltop_254_284 top254 top284 {l}
Rbot_254_284 bot254 bot284 {r}
Lbot_254_284 bot254 bot284 {l}
C254 top254 bot254 {c}
Rtop_255_256 top255 top256 {r}
Ltop_255_256 top255 top256 {l}
Rbot_255_256 bot255 bot256 {r}
Lbot_255_256 bot255 bot256 {l}
Rtop_255_285 top255 top285 {r}
Ltop_255_285 top255 top285 {l}
Rbot_255_285 bot255 bot285 {r}
Lbot_255_285 bot255 bot285 {l}
C255 top255 bot255 {c}
Rtop_256_257 top256 top257 {r}
Ltop_256_257 top256 top257 {l}
Rbot_256_257 bot256 bot257 {r}
Lbot_256_257 bot256 bot257 {l}
Rtop_256_286 top256 top286 {r}
Ltop_256_286 top256 top286 {l}
Rbot_256_286 bot256 bot286 {r}
Lbot_256_286 bot256 bot286 {l}
C256 top256 bot256 {c}
Rtop_257_258 top257 top258 {r}
Ltop_257_258 top257 top258 {l}
Rbot_257_258 bot257 bot258 {r}
Lbot_257_258 bot257 bot258 {l}
Rtop_257_287 top257 top287 {r}
Ltop_257_287 top257 top287 {l}
Rbot_257_287 bot257 bot287 {r}
Lbot_257_287 bot257 bot287 {l}
C257 top257 bot257 {c}
Rtop_258_259 top258 top259 {r}
Ltop_258_259 top258 top259 {l}
Rbot_258_259 bot258 bot259 {r}
Lbot_258_259 bot258 bot259 {l}
Rtop_258_288 top258 top288 {r}
Ltop_258_288 top258 top288 {l}
Rbot_258_288 bot258 bot288 {r}
Lbot_258_288 bot258 bot288 {l}
C258 top258 bot258 {c}
Rtop_259_260 top259 top260 {r}
Ltop_259_260 top259 top260 {l}
Rbot_259_260 bot259 bot260 {r}
Lbot_259_260 bot259 bot260 {l}
Rtop_259_289 top259 top289 {r}
Ltop_259_289 top259 top289 {l}
Rbot_259_289 bot259 bot289 {r}
Lbot_259_289 bot259 bot289 {l}
C259 top259 bot259 {c}
Rtop_260_261 top260 top261 {r}
Ltop_260_261 top260 top261 {l}
Rbot_260_261 bot260 bot261 {r}
Lbot_260_261 bot260 bot261 {l}
Rtop_260_290 top260 top290 {r}
Ltop_260_290 top260 top290 {l}
Rbot_260_290 bot260 bot290 {r}
Lbot_260_290 bot260 bot290 {l}
C260 top260 bot260 {c}
Rtop_261_262 top261 top262 {r}
Ltop_261_262 top261 top262 {l}
Rbot_261_262 bot261 bot262 {r}
Lbot_261_262 bot261 bot262 {l}
Rtop_261_291 top261 top291 {r}
Ltop_261_291 top261 top291 {l}
Rbot_261_291 bot261 bot291 {r}
Lbot_261_291 bot261 bot291 {l}
C261 top261 bot261 {c}
Rtop_262_263 top262 top263 {r}
Ltop_262_263 top262 top263 {l}
Rbot_262_263 bot262 bot263 {r}
Lbot_262_263 bot262 bot263 {l}
Rtop_262_292 top262 top292 {r}
Ltop_262_292 top262 top292 {l}
Rbot_262_292 bot262 bot292 {r}
Lbot_262_292 bot262 bot292 {l}
C262 top262 bot262 {c}
Rtop_263_264 top263 top264 {r}
Ltop_263_264 top263 top264 {l}
Rbot_263_264 bot263 bot264 {r}
Lbot_263_264 bot263 bot264 {l}
Rtop_263_293 top263 top293 {r}
Ltop_263_293 top263 top293 {l}
Rbot_263_293 bot263 bot293 {r}
Lbot_263_293 bot263 bot293 {l}
C263 top263 bot263 {c}
Rtop_264_265 top264 top265 {r}
Ltop_264_265 top264 top265 {l}
Rbot_264_265 bot264 bot265 {r}
Lbot_264_265 bot264 bot265 {l}
Rtop_264_294 top264 top294 {r}
Ltop_264_294 top264 top294 {l}
Rbot_264_294 bot264 bot294 {r}
Lbot_264_294 bot264 bot294 {l}
C264 top264 bot264 {c}
Rtop_265_266 top265 top266 {r}
Ltop_265_266 top265 top266 {l}
Rbot_265_266 bot265 bot266 {r}
Lbot_265_266 bot265 bot266 {l}
Rtop_265_295 top265 top295 {r}
Ltop_265_295 top265 top295 {l}
Rbot_265_295 bot265 bot295 {r}
Lbot_265_295 bot265 bot295 {l}
C265 top265 bot265 {c}
Rtop_266_267 top266 top267 {r}
Ltop_266_267 top266 top267 {l}
Rbot_266_267 bot266 bot267 {r}
Lbot_266_267 bot266 bot267 {l}
Rtop_266_296 top266 top296 {r}
Ltop_266_296 top266 top296 {l}
Rbot_266_296 bot266 bot296 {r}
Lbot_266_296 bot266 bot296 {l}
C266 top266 bot266 {c}
Rtop_267_268 top267 top268 {r}
Ltop_267_268 top267 top268 {l}
Rbot_267_268 bot267 bot268 {r}
Lbot_267_268 bot267 bot268 {l}
Rtop_267_297 top267 top297 {r}
Ltop_267_297 top267 top297 {l}
Rbot_267_297 bot267 bot297 {r}
Lbot_267_297 bot267 bot297 {l}
C267 top267 bot267 {c}
Rtop_268_269 top268 top269 {r}
Ltop_268_269 top268 top269 {l}
Rbot_268_269 bot268 bot269 {r}
Lbot_268_269 bot268 bot269 {l}
Rtop_268_298 top268 top298 {r}
Ltop_268_298 top268 top298 {l}
Rbot_268_298 bot268 bot298 {r}
Lbot_268_298 bot268 bot298 {l}
C268 top268 bot268 {c}
Rtop_269_270 top269 top270 {r}
Ltop_269_270 top269 top270 {l}
Rbot_269_270 bot269 bot270 {r}
Lbot_269_270 bot269 bot270 {l}
Rtop_269_299 top269 top299 {r}
Ltop_269_299 top269 top299 {l}
Rbot_269_299 bot269 bot299 {r}
Lbot_269_299 bot269 bot299 {l}
C269 top269 bot269 {c}
Rtop_270_300 top270 top300 {r}
Ltop_270_300 top270 top300 {l}
Rbot_270_300 bot270 bot300 {r}
Lbot_270_300 bot270 bot300 {l}
C270 top270 bot270 {c}
Rtop_271_272 top271 top272 {r}
Ltop_271_272 top271 top272 {l}
Rbot_271_272 bot271 bot272 {r}
Lbot_271_272 bot271 bot272 {l}
Rtop_271_301 top271 top301 {r}
Ltop_271_301 top271 top301 {l}
Rbot_271_301 bot271 bot301 {r}
Lbot_271_301 bot271 bot301 {l}
C271 top271 bot271 {c}
Rtop_272_273 top272 top273 {r}
Ltop_272_273 top272 top273 {l}
Rbot_272_273 bot272 bot273 {r}
Lbot_272_273 bot272 bot273 {l}
Rtop_272_302 top272 top302 {r}
Ltop_272_302 top272 top302 {l}
Rbot_272_302 bot272 bot302 {r}
Lbot_272_302 bot272 bot302 {l}
C272 top272 bot272 {c}
Rtop_273_274 top273 top274 {r}
Ltop_273_274 top273 top274 {l}
Rbot_273_274 bot273 bot274 {r}
Lbot_273_274 bot273 bot274 {l}
Rtop_273_303 top273 top303 {r}
Ltop_273_303 top273 top303 {l}
Rbot_273_303 bot273 bot303 {r}
Lbot_273_303 bot273 bot303 {l}
C273 top273 bot273 {c}
Rtop_274_275 top274 top275 {r}
Ltop_274_275 top274 top275 {l}
Rbot_274_275 bot274 bot275 {r}
Lbot_274_275 bot274 bot275 {l}
Rtop_274_304 top274 top304 {r}
Ltop_274_304 top274 top304 {l}
Rbot_274_304 bot274 bot304 {r}
Lbot_274_304 bot274 bot304 {l}
C274 top274 bot274 {c}
Rtop_275_276 top275 top276 {r}
Ltop_275_276 top275 top276 {l}
Rbot_275_276 bot275 bot276 {r}
Lbot_275_276 bot275 bot276 {l}
Rtop_275_305 top275 top305 {r}
Ltop_275_305 top275 top305 {l}
Rbot_275_305 bot275 bot305 {r}
Lbot_275_305 bot275 bot305 {l}
C275 top275 bot275 {c}
Rtop_276_277 top276 top277 {r}
Ltop_276_277 top276 top277 {l}
Rbot_276_277 bot276 bot277 {r}
Lbot_276_277 bot276 bot277 {l}
Rtop_276_306 top276 top306 {r}
Ltop_276_306 top276 top306 {l}
Rbot_276_306 bot276 bot306 {r}
Lbot_276_306 bot276 bot306 {l}
C276 top276 bot276 {c}
Rtop_277_278 top277 top278 {r}
Ltop_277_278 top277 top278 {l}
Rbot_277_278 bot277 bot278 {r}
Lbot_277_278 bot277 bot278 {l}
Rtop_277_307 top277 top307 {r}
Ltop_277_307 top277 top307 {l}
Rbot_277_307 bot277 bot307 {r}
Lbot_277_307 bot277 bot307 {l}
C277 top277 bot277 {c}
Rtop_278_279 top278 top279 {r}
Ltop_278_279 top278 top279 {l}
Rbot_278_279 bot278 bot279 {r}
Lbot_278_279 bot278 bot279 {l}
Rtop_278_308 top278 top308 {r}
Ltop_278_308 top278 top308 {l}
Rbot_278_308 bot278 bot308 {r}
Lbot_278_308 bot278 bot308 {l}
C278 top278 bot278 {c}
Rtop_279_280 top279 top280 {r}
Ltop_279_280 top279 top280 {l}
Rbot_279_280 bot279 bot280 {r}
Lbot_279_280 bot279 bot280 {l}
Rtop_279_309 top279 top309 {r}
Ltop_279_309 top279 top309 {l}
Rbot_279_309 bot279 bot309 {r}
Lbot_279_309 bot279 bot309 {l}
C279 top279 bot279 {c}
Rtop_280_281 top280 top281 {r}
Ltop_280_281 top280 top281 {l}
Rbot_280_281 bot280 bot281 {r}
Lbot_280_281 bot280 bot281 {l}
Rtop_280_310 top280 top310 {r}
Ltop_280_310 top280 top310 {l}
Rbot_280_310 bot280 bot310 {r}
Lbot_280_310 bot280 bot310 {l}
C280 top280 bot280 {c}
Rtop_281_282 top281 top282 {r}
Ltop_281_282 top281 top282 {l}
Rbot_281_282 bot281 bot282 {r}
Lbot_281_282 bot281 bot282 {l}
Rtop_281_311 top281 top311 {r}
Ltop_281_311 top281 top311 {l}
Rbot_281_311 bot281 bot311 {r}
Lbot_281_311 bot281 bot311 {l}
C281 top281 bot281 {c}
Rtop_282_283 top282 top283 {r}
Ltop_282_283 top282 top283 {l}
Rbot_282_283 bot282 bot283 {r}
Lbot_282_283 bot282 bot283 {l}
Rtop_282_312 top282 top312 {r}
Ltop_282_312 top282 top312 {l}
Rbot_282_312 bot282 bot312 {r}
Lbot_282_312 bot282 bot312 {l}
C282 top282 bot282 {c}
Rtop_283_284 top283 top284 {r}
Ltop_283_284 top283 top284 {l}
Rbot_283_284 bot283 bot284 {r}
Lbot_283_284 bot283 bot284 {l}
Rtop_283_313 top283 top313 {r}
Ltop_283_313 top283 top313 {l}
Rbot_283_313 bot283 bot313 {r}
Lbot_283_313 bot283 bot313 {l}
C283 top283 bot283 {c}
Rtop_284_285 top284 top285 {r}
Ltop_284_285 top284 top285 {l}
Rbot_284_285 bot284 bot285 {r}
Lbot_284_285 bot284 bot285 {l}
Rtop_284_314 top284 top314 {r}
Ltop_284_314 top284 top314 {l}
Rbot_284_314 bot284 bot314 {r}
Lbot_284_314 bot284 bot314 {l}
C284 top284 bot284 {c}
Rtop_285_286 top285 top286 {r}
Ltop_285_286 top285 top286 {l}
Rbot_285_286 bot285 bot286 {r}
Lbot_285_286 bot285 bot286 {l}
Rtop_285_315 top285 top315 {r}
Ltop_285_315 top285 top315 {l}
Rbot_285_315 bot285 bot315 {r}
Lbot_285_315 bot285 bot315 {l}
C285 top285 bot285 {c}
Rtop_286_287 top286 top287 {r}
Ltop_286_287 top286 top287 {l}
Rbot_286_287 bot286 bot287 {r}
Lbot_286_287 bot286 bot287 {l}
Rtop_286_316 top286 top316 {r}
Ltop_286_316 top286 top316 {l}
Rbot_286_316 bot286 bot316 {r}
Lbot_286_316 bot286 bot316 {l}
C286 top286 bot286 {c}
Rtop_287_288 top287 top288 {r}
Ltop_287_288 top287 top288 {l}
Rbot_287_288 bot287 bot288 {r}
Lbot_287_288 bot287 bot288 {l}
Rtop_287_317 top287 top317 {r}
Ltop_287_317 top287 top317 {l}
Rbot_287_317 bot287 bot317 {r}
Lbot_287_317 bot287 bot317 {l}
C287 top287 bot287 {c}
Rtop_288_289 top288 top289 {r}
Ltop_288_289 top288 top289 {l}
Rbot_288_289 bot288 bot289 {r}
Lbot_288_289 bot288 bot289 {l}
Rtop_288_318 top288 top318 {r}
Ltop_288_318 top288 top318 {l}
Rbot_288_318 bot288 bot318 {r}
Lbot_288_318 bot288 bot318 {l}
C288 top288 bot288 {c}
Rtop_289_290 top289 top290 {r}
Ltop_289_290 top289 top290 {l}
Rbot_289_290 bot289 bot290 {r}
Lbot_289_290 bot289 bot290 {l}
Rtop_289_319 top289 top319 {r}
Ltop_289_319 top289 top319 {l}
Rbot_289_319 bot289 bot319 {r}
Lbot_289_319 bot289 bot319 {l}
C289 top289 bot289 {c}
Rtop_290_291 top290 top291 {r}
Ltop_290_291 top290 top291 {l}
Rbot_290_291 bot290 bot291 {r}
Lbot_290_291 bot290 bot291 {l}
Rtop_290_320 top290 top320 {r}
Ltop_290_320 top290 top320 {l}
Rbot_290_320 bot290 bot320 {r}
Lbot_290_320 bot290 bot320 {l}
C290 top290 bot290 {c}
Rtop_291_292 top291 top292 {r}
Ltop_291_292 top291 top292 {l}
Rbot_291_292 bot291 bot292 {r}
Lbot_291_292 bot291 bot292 {l}
Rtop_291_321 top291 top321 {r}
Ltop_291_321 top291 top321 {l}
Rbot_291_321 bot291 bot321 {r}
Lbot_291_321 bot291 bot321 {l}
C291 top291 bot291 {c}
Rtop_292_293 top292 top293 {r}
Ltop_292_293 top292 top293 {l}
Rbot_292_293 bot292 bot293 {r}
Lbot_292_293 bot292 bot293 {l}
Rtop_292_322 top292 top322 {r}
Ltop_292_322 top292 top322 {l}
Rbot_292_322 bot292 bot322 {r}
Lbot_292_322 bot292 bot322 {l}
C292 top292 bot292 {c}
Rtop_293_294 top293 top294 {r}
Ltop_293_294 top293 top294 {l}
Rbot_293_294 bot293 bot294 {r}
Lbot_293_294 bot293 bot294 {l}
Rtop_293_323 top293 top323 {r}
Ltop_293_323 top293 top323 {l}
Rbot_293_323 bot293 bot323 {r}
Lbot_293_323 bot293 bot323 {l}
C293 top293 bot293 {c}
Rtop_294_295 top294 top295 {r}
Ltop_294_295 top294 top295 {l}
Rbot_294_295 bot294 bot295 {r}
Lbot_294_295 bot294 bot295 {l}
Rtop_294_324 top294 top324 {r}
Ltop_294_324 top294 top324 {l}
Rbot_294_324 bot294 bot324 {r}
Lbot_294_324 bot294 bot324 {l}
C294 top294 bot294 {c}
Rtop_295_296 top295 top296 {r}
Ltop_295_296 top295 top296 {l}
Rbot_295_296 bot295 bot296 {r}
Lbot_295_296 bot295 bot296 {l}
Rtop_295_325 top295 top325 {r}
Ltop_295_325 top295 top325 {l}
Rbot_295_325 bot295 bot325 {r}
Lbot_295_325 bot295 bot325 {l}
C295 top295 bot295 {c}
Rtop_296_297 top296 top297 {r}
Ltop_296_297 top296 top297 {l}
Rbot_296_297 bot296 bot297 {r}
Lbot_296_297 bot296 bot297 {l}
Rtop_296_326 top296 top326 {r}
Ltop_296_326 top296 top326 {l}
Rbot_296_326 bot296 bot326 {r}
Lbot_296_326 bot296 bot326 {l}
C296 top296 bot296 {c}
Rtop_297_298 top297 top298 {r}
Ltop_297_298 top297 top298 {l}
Rbot_297_298 bot297 bot298 {r}
Lbot_297_298 bot297 bot298 {l}
Rtop_297_327 top297 top327 {r}
Ltop_297_327 top297 top327 {l}
Rbot_297_327 bot297 bot327 {r}
Lbot_297_327 bot297 bot327 {l}
C297 top297 bot297 {c}
Rtop_298_299 top298 top299 {r}
Ltop_298_299 top298 top299 {l}
Rbot_298_299 bot298 bot299 {r}
Lbot_298_299 bot298 bot299 {l}
Rtop_298_328 top298 top328 {r}
Ltop_298_328 top298 top328 {l}
Rbot_298_328 bot298 bot328 {r}
Lbot_298_328 bot298 bot328 {l}
C298 top298 bot298 {c}
Rtop_299_300 top299 top300 {r}
Ltop_299_300 top299 top300 {l}
Rbot_299_300 bot299 bot300 {r}
Lbot_299_300 bot299 bot300 {l}
Rtop_299_329 top299 top329 {r}
Ltop_299_329 top299 top329 {l}
Rbot_299_329 bot299 bot329 {r}
Lbot_299_329 bot299 bot329 {l}
C299 top299 bot299 {c}
Rtop_300_330 top300 top330 {r}
Ltop_300_330 top300 top330 {l}
Rbot_300_330 bot300 bot330 {r}
Lbot_300_330 bot300 bot330 {l}
C300 top300 bot300 {c}
Rtop_301_302 top301 top302 {r}
Ltop_301_302 top301 top302 {l}
Rbot_301_302 bot301 bot302 {r}
Lbot_301_302 bot301 bot302 {l}
Rtop_301_331 top301 top331 {r}
Ltop_301_331 top301 top331 {l}
Rbot_301_331 bot301 bot331 {r}
Lbot_301_331 bot301 bot331 {l}
C301 top301 bot301 {c}
Rtop_302_303 top302 top303 {r}
Ltop_302_303 top302 top303 {l}
Rbot_302_303 bot302 bot303 {r}
Lbot_302_303 bot302 bot303 {l}
Rtop_302_332 top302 top332 {r}
Ltop_302_332 top302 top332 {l}
Rbot_302_332 bot302 bot332 {r}
Lbot_302_332 bot302 bot332 {l}
C302 top302 bot302 {c}
Rtop_303_304 top303 top304 {r}
Ltop_303_304 top303 top304 {l}
Rbot_303_304 bot303 bot304 {r}
Lbot_303_304 bot303 bot304 {l}
Rtop_303_333 top303 top333 {r}
Ltop_303_333 top303 top333 {l}
Rbot_303_333 bot303 bot333 {r}
Lbot_303_333 bot303 bot333 {l}
C303 top303 bot303 {c}
Rtop_304_305 top304 top305 {r}
Ltop_304_305 top304 top305 {l}
Rbot_304_305 bot304 bot305 {r}
Lbot_304_305 bot304 bot305 {l}
Rtop_304_334 top304 top334 {r}
Ltop_304_334 top304 top334 {l}
Rbot_304_334 bot304 bot334 {r}
Lbot_304_334 bot304 bot334 {l}
C304 top304 bot304 {c}
Rtop_305_306 top305 top306 {r}
Ltop_305_306 top305 top306 {l}
Rbot_305_306 bot305 bot306 {r}
Lbot_305_306 bot305 bot306 {l}
Rtop_305_335 top305 top335 {r}
Ltop_305_335 top305 top335 {l}
Rbot_305_335 bot305 bot335 {r}
Lbot_305_335 bot305 bot335 {l}
C305 top305 bot305 {c}
Rtop_306_307 top306 top307 {r}
Ltop_306_307 top306 top307 {l}
Rbot_306_307 bot306 bot307 {r}
Lbot_306_307 bot306 bot307 {l}
Rtop_306_336 top306 top336 {r}
Ltop_306_336 top306 top336 {l}
Rbot_306_336 bot306 bot336 {r}
Lbot_306_336 bot306 bot336 {l}
C306 top306 bot306 {c}
Rtop_307_308 top307 top308 {r}
Ltop_307_308 top307 top308 {l}
Rbot_307_308 bot307 bot308 {r}
Lbot_307_308 bot307 bot308 {l}
Rtop_307_337 top307 top337 {r}
Ltop_307_337 top307 top337 {l}
Rbot_307_337 bot307 bot337 {r}
Lbot_307_337 bot307 bot337 {l}
C307 top307 bot307 {c}
Rtop_308_309 top308 top309 {r}
Ltop_308_309 top308 top309 {l}
Rbot_308_309 bot308 bot309 {r}
Lbot_308_309 bot308 bot309 {l}
Rtop_308_338 top308 top338 {r}
Ltop_308_338 top308 top338 {l}
Rbot_308_338 bot308 bot338 {r}
Lbot_308_338 bot308 bot338 {l}
C308 top308 bot308 {c}
Rtop_309_310 top309 top310 {r}
Ltop_309_310 top309 top310 {l}
Rbot_309_310 bot309 bot310 {r}
Lbot_309_310 bot309 bot310 {l}
Rtop_309_339 top309 top339 {r}
Ltop_309_339 top309 top339 {l}
Rbot_309_339 bot309 bot339 {r}
Lbot_309_339 bot309 bot339 {l}
C309 top309 bot309 {c}
Rtop_310_311 top310 top311 {r}
Ltop_310_311 top310 top311 {l}
Rbot_310_311 bot310 bot311 {r}
Lbot_310_311 bot310 bot311 {l}
Rtop_310_340 top310 top340 {r}
Ltop_310_340 top310 top340 {l}
Rbot_310_340 bot310 bot340 {r}
Lbot_310_340 bot310 bot340 {l}
C310 top310 bot310 {c}
Rtop_311_312 top311 top312 {r}
Ltop_311_312 top311 top312 {l}
Rbot_311_312 bot311 bot312 {r}
Lbot_311_312 bot311 bot312 {l}
Rtop_311_341 top311 top341 {r}
Ltop_311_341 top311 top341 {l}
Rbot_311_341 bot311 bot341 {r}
Lbot_311_341 bot311 bot341 {l}
C311 top311 bot311 {c}
Rtop_312_313 top312 top313 {r}
Ltop_312_313 top312 top313 {l}
Rbot_312_313 bot312 bot313 {r}
Lbot_312_313 bot312 bot313 {l}
Rtop_312_342 top312 top342 {r}
Ltop_312_342 top312 top342 {l}
Rbot_312_342 bot312 bot342 {r}
Lbot_312_342 bot312 bot342 {l}
C312 top312 bot312 {c}
Rtop_313_314 top313 top314 {r}
Ltop_313_314 top313 top314 {l}
Rbot_313_314 bot313 bot314 {r}
Lbot_313_314 bot313 bot314 {l}
Rtop_313_343 top313 top343 {r}
Ltop_313_343 top313 top343 {l}
Rbot_313_343 bot313 bot343 {r}
Lbot_313_343 bot313 bot343 {l}
C313 top313 bot313 {c}
Rtop_314_315 top314 top315 {r}
Ltop_314_315 top314 top315 {l}
Rbot_314_315 bot314 bot315 {r}
Lbot_314_315 bot314 bot315 {l}
Rtop_314_344 top314 top344 {r}
Ltop_314_344 top314 top344 {l}
Rbot_314_344 bot314 bot344 {r}
Lbot_314_344 bot314 bot344 {l}
C314 top314 bot314 {c}
Rtop_315_316 top315 top316 {r}
Ltop_315_316 top315 top316 {l}
Rbot_315_316 bot315 bot316 {r}
Lbot_315_316 bot315 bot316 {l}
Rtop_315_345 top315 top345 {r}
Ltop_315_345 top315 top345 {l}
Rbot_315_345 bot315 bot345 {r}
Lbot_315_345 bot315 bot345 {l}
C315 top315 bot315 {c}
Rtop_316_317 top316 top317 {r}
Ltop_316_317 top316 top317 {l}
Rbot_316_317 bot316 bot317 {r}
Lbot_316_317 bot316 bot317 {l}
Rtop_316_346 top316 top346 {r}
Ltop_316_346 top316 top346 {l}
Rbot_316_346 bot316 bot346 {r}
Lbot_316_346 bot316 bot346 {l}
C316 top316 bot316 {c}
Rtop_317_318 top317 top318 {r}
Ltop_317_318 top317 top318 {l}
Rbot_317_318 bot317 bot318 {r}
Lbot_317_318 bot317 bot318 {l}
Rtop_317_347 top317 top347 {r}
Ltop_317_347 top317 top347 {l}
Rbot_317_347 bot317 bot347 {r}
Lbot_317_347 bot317 bot347 {l}
C317 top317 bot317 {c}
Rtop_318_319 top318 top319 {r}
Ltop_318_319 top318 top319 {l}
Rbot_318_319 bot318 bot319 {r}
Lbot_318_319 bot318 bot319 {l}
Rtop_318_348 top318 top348 {r}
Ltop_318_348 top318 top348 {l}
Rbot_318_348 bot318 bot348 {r}
Lbot_318_348 bot318 bot348 {l}
C318 top318 bot318 {c}
Rtop_319_320 top319 top320 {r}
Ltop_319_320 top319 top320 {l}
Rbot_319_320 bot319 bot320 {r}
Lbot_319_320 bot319 bot320 {l}
Rtop_319_349 top319 top349 {r}
Ltop_319_349 top319 top349 {l}
Rbot_319_349 bot319 bot349 {r}
Lbot_319_349 bot319 bot349 {l}
C319 top319 bot319 {c}
Rtop_320_321 top320 top321 {r}
Ltop_320_321 top320 top321 {l}
Rbot_320_321 bot320 bot321 {r}
Lbot_320_321 bot320 bot321 {l}
Rtop_320_350 top320 top350 {r}
Ltop_320_350 top320 top350 {l}
Rbot_320_350 bot320 bot350 {r}
Lbot_320_350 bot320 bot350 {l}
C320 top320 bot320 {c}
Rtop_321_322 top321 top322 {r}
Ltop_321_322 top321 top322 {l}
Rbot_321_322 bot321 bot322 {r}
Lbot_321_322 bot321 bot322 {l}
Rtop_321_351 top321 top351 {r}
Ltop_321_351 top321 top351 {l}
Rbot_321_351 bot321 bot351 {r}
Lbot_321_351 bot321 bot351 {l}
C321 top321 bot321 {c}
Rtop_322_323 top322 top323 {r}
Ltop_322_323 top322 top323 {l}
Rbot_322_323 bot322 bot323 {r}
Lbot_322_323 bot322 bot323 {l}
Rtop_322_352 top322 top352 {r}
Ltop_322_352 top322 top352 {l}
Rbot_322_352 bot322 bot352 {r}
Lbot_322_352 bot322 bot352 {l}
C322 top322 bot322 {c}
Rtop_323_324 top323 top324 {r}
Ltop_323_324 top323 top324 {l}
Rbot_323_324 bot323 bot324 {r}
Lbot_323_324 bot323 bot324 {l}
Rtop_323_353 top323 top353 {r}
Ltop_323_353 top323 top353 {l}
Rbot_323_353 bot323 bot353 {r}
Lbot_323_353 bot323 bot353 {l}
C323 top323 bot323 {c}
Rtop_324_325 top324 top325 {r}
Ltop_324_325 top324 top325 {l}
Rbot_324_325 bot324 bot325 {r}
Lbot_324_325 bot324 bot325 {l}
Rtop_324_354 top324 top354 {r}
Ltop_324_354 top324 top354 {l}
Rbot_324_354 bot324 bot354 {r}
Lbot_324_354 bot324 bot354 {l}
C324 top324 bot324 {c}
Rtop_325_326 top325 top326 {r}
Ltop_325_326 top325 top326 {l}
Rbot_325_326 bot325 bot326 {r}
Lbot_325_326 bot325 bot326 {l}
Rtop_325_355 top325 top355 {r}
Ltop_325_355 top325 top355 {l}
Rbot_325_355 bot325 bot355 {r}
Lbot_325_355 bot325 bot355 {l}
C325 top325 bot325 {c}
Rtop_326_327 top326 top327 {r}
Ltop_326_327 top326 top327 {l}
Rbot_326_327 bot326 bot327 {r}
Lbot_326_327 bot326 bot327 {l}
Rtop_326_356 top326 top356 {r}
Ltop_326_356 top326 top356 {l}
Rbot_326_356 bot326 bot356 {r}
Lbot_326_356 bot326 bot356 {l}
C326 top326 bot326 {c}
Rtop_327_328 top327 top328 {r}
Ltop_327_328 top327 top328 {l}
Rbot_327_328 bot327 bot328 {r}
Lbot_327_328 bot327 bot328 {l}
Rtop_327_357 top327 top357 {r}
Ltop_327_357 top327 top357 {l}
Rbot_327_357 bot327 bot357 {r}
Lbot_327_357 bot327 bot357 {l}
C327 top327 bot327 {c}
Rtop_328_329 top328 top329 {r}
Ltop_328_329 top328 top329 {l}
Rbot_328_329 bot328 bot329 {r}
Lbot_328_329 bot328 bot329 {l}
Rtop_328_358 top328 top358 {r}
Ltop_328_358 top328 top358 {l}
Rbot_328_358 bot328 bot358 {r}
Lbot_328_358 bot328 bot358 {l}
C328 top328 bot328 {c}
Rtop_329_330 top329 top330 {r}
Ltop_329_330 top329 top330 {l}
Rbot_329_330 bot329 bot330 {r}
Lbot_329_330 bot329 bot330 {l}
Rtop_329_359 top329 top359 {r}
Ltop_329_359 top329 top359 {l}
Rbot_329_359 bot329 bot359 {r}
Lbot_329_359 bot329 bot359 {l}
C329 top329 bot329 {c}
Rtop_330_360 top330 top360 {r}
Ltop_330_360 top330 top360 {l}
Rbot_330_360 bot330 bot360 {r}
Lbot_330_360 bot330 bot360 {l}
C330 top330 bot330 {c}
Rtop_331_332 top331 top332 {r}
Ltop_331_332 top331 top332 {l}
Rbot_331_332 bot331 bot332 {r}
Lbot_331_332 bot331 bot332 {l}
Rtop_331_361 top331 top361 {r}
Ltop_331_361 top331 top361 {l}
Rbot_331_361 bot331 bot361 {r}
Lbot_331_361 bot331 bot361 {l}
C331 top331 bot331 {c}
Rtop_332_333 top332 top333 {r}
Ltop_332_333 top332 top333 {l}
Rbot_332_333 bot332 bot333 {r}
Lbot_332_333 bot332 bot333 {l}
Rtop_332_362 top332 top362 {r}
Ltop_332_362 top332 top362 {l}
Rbot_332_362 bot332 bot362 {r}
Lbot_332_362 bot332 bot362 {l}
C332 top332 bot332 {c}
Rtop_333_334 top333 top334 {r}
Ltop_333_334 top333 top334 {l}
Rbot_333_334 bot333 bot334 {r}
Lbot_333_334 bot333 bot334 {l}
Rtop_333_363 top333 top363 {r}
Ltop_333_363 top333 top363 {l}
Rbot_333_363 bot333 bot363 {r}
Lbot_333_363 bot333 bot363 {l}
C333 top333 bot333 {c}
Rtop_334_335 top334 top335 {r}
Ltop_334_335 top334 top335 {l}
Rbot_334_335 bot334 bot335 {r}
Lbot_334_335 bot334 bot335 {l}
Rtop_334_364 top334 top364 {r}
Ltop_334_364 top334 top364 {l}
Rbot_334_364 bot334 bot364 {r}
Lbot_334_364 bot334 bot364 {l}
C334 top334 bot334 {c}
Rtop_335_336 top335 top336 {r}
Ltop_335_336 top335 top336 {l}
Rbot_335_336 bot335 bot336 {r}
Lbot_335_336 bot335 bot336 {l}
Rtop_335_365 top335 top365 {r}
Ltop_335_365 top335 top365 {l}
Rbot_335_365 bot335 bot365 {r}
Lbot_335_365 bot335 bot365 {l}
C335 top335 bot335 {c}
Rtop_336_337 top336 top337 {r}
Ltop_336_337 top336 top337 {l}
Rbot_336_337 bot336 bot337 {r}
Lbot_336_337 bot336 bot337 {l}
Rtop_336_366 top336 top366 {r}
Ltop_336_366 top336 top366 {l}
Rbot_336_366 bot336 bot366 {r}
Lbot_336_366 bot336 bot366 {l}
C336 top336 bot336 {c}
Rtop_337_338 top337 top338 {r}
Ltop_337_338 top337 top338 {l}
Rbot_337_338 bot337 bot338 {r}
Lbot_337_338 bot337 bot338 {l}
Rtop_337_367 top337 top367 {r}
Ltop_337_367 top337 top367 {l}
Rbot_337_367 bot337 bot367 {r}
Lbot_337_367 bot337 bot367 {l}
C337 top337 bot337 {c}
Rtop_338_339 top338 top339 {r}
Ltop_338_339 top338 top339 {l}
Rbot_338_339 bot338 bot339 {r}
Lbot_338_339 bot338 bot339 {l}
Rtop_338_368 top338 top368 {r}
Ltop_338_368 top338 top368 {l}
Rbot_338_368 bot338 bot368 {r}
Lbot_338_368 bot338 bot368 {l}
C338 top338 bot338 {c}
Rtop_339_340 top339 top340 {r}
Ltop_339_340 top339 top340 {l}
Rbot_339_340 bot339 bot340 {r}
Lbot_339_340 bot339 bot340 {l}
Rtop_339_369 top339 top369 {r}
Ltop_339_369 top339 top369 {l}
Rbot_339_369 bot339 bot369 {r}
Lbot_339_369 bot339 bot369 {l}
C339 top339 bot339 {c}
Rtop_340_341 top340 top341 {r}
Ltop_340_341 top340 top341 {l}
Rbot_340_341 bot340 bot341 {r}
Lbot_340_341 bot340 bot341 {l}
Rtop_340_370 top340 top370 {r}
Ltop_340_370 top340 top370 {l}
Rbot_340_370 bot340 bot370 {r}
Lbot_340_370 bot340 bot370 {l}
C340 top340 bot340 {c}
Rtop_341_342 top341 top342 {r}
Ltop_341_342 top341 top342 {l}
Rbot_341_342 bot341 bot342 {r}
Lbot_341_342 bot341 bot342 {l}
Rtop_341_371 top341 top371 {r}
Ltop_341_371 top341 top371 {l}
Rbot_341_371 bot341 bot371 {r}
Lbot_341_371 bot341 bot371 {l}
C341 top341 bot341 {c}
Rtop_342_343 top342 top343 {r}
Ltop_342_343 top342 top343 {l}
Rbot_342_343 bot342 bot343 {r}
Lbot_342_343 bot342 bot343 {l}
Rtop_342_372 top342 top372 {r}
Ltop_342_372 top342 top372 {l}
Rbot_342_372 bot342 bot372 {r}
Lbot_342_372 bot342 bot372 {l}
C342 top342 bot342 {c}
Rtop_343_344 top343 top344 {r}
Ltop_343_344 top343 top344 {l}
Rbot_343_344 bot343 bot344 {r}
Lbot_343_344 bot343 bot344 {l}
Rtop_343_373 top343 top373 {r}
Ltop_343_373 top343 top373 {l}
Rbot_343_373 bot343 bot373 {r}
Lbot_343_373 bot343 bot373 {l}
C343 top343 bot343 {c}
Rtop_344_345 top344 top345 {r}
Ltop_344_345 top344 top345 {l}
Rbot_344_345 bot344 bot345 {r}
Lbot_344_345 bot344 bot345 {l}
Rtop_344_374 top344 top374 {r}
Ltop_344_374 top344 top374 {l}
Rbot_344_374 bot344 bot374 {r}
Lbot_344_374 bot344 bot374 {l}
C344 top344 bot344 {c}
Rtop_345_346 top345 top346 {r}
Ltop_345_346 top345 top346 {l}
Rbot_345_346 bot345 bot346 {r}
Lbot_345_346 bot345 bot346 {l}
Rtop_345_375 top345 top375 {r}
Ltop_345_375 top345 top375 {l}
Rbot_345_375 bot345 bot375 {r}
Lbot_345_375 bot345 bot375 {l}
C345 top345 bot345 {c}
Rtop_346_347 top346 top347 {r}
Ltop_346_347 top346 top347 {l}
Rbot_346_347 bot346 bot347 {r}
Lbot_346_347 bot346 bot347 {l}
Rtop_346_376 top346 top376 {r}
Ltop_346_376 top346 top376 {l}
Rbot_346_376 bot346 bot376 {r}
Lbot_346_376 bot346 bot376 {l}
C346 top346 bot346 {c}
Rtop_347_348 top347 top348 {r}
Ltop_347_348 top347 top348 {l}
Rbot_347_348 bot347 bot348 {r}
Lbot_347_348 bot347 bot348 {l}
Rtop_347_377 top347 top377 {r}
Ltop_347_377 top347 top377 {l}
Rbot_347_377 bot347 bot377 {r}
Lbot_347_377 bot347 bot377 {l}
C347 top347 bot347 {c}
Rtop_348_349 top348 top349 {r}
Ltop_348_349 top348 top349 {l}
Rbot_348_349 bot348 bot349 {r}
Lbot_348_349 bot348 bot349 {l}
Rtop_348_378 top348 top378 {r}
Ltop_348_378 top348 top378 {l}
Rbot_348_378 bot348 bot378 {r}
Lbot_348_378 bot348 bot378 {l}
C348 top348 bot348 {c}
Rtop_349_350 top349 top350 {r}
Ltop_349_350 top349 top350 {l}
Rbot_349_350 bot349 bot350 {r}
Lbot_349_350 bot349 bot350 {l}
Rtop_349_379 top349 top379 {r}
Ltop_349_379 top349 top379 {l}
Rbot_349_379 bot349 bot379 {r}
Lbot_349_379 bot349 bot379 {l}
C349 top349 bot349 {c}
Rtop_350_351 top350 top351 {r}
Ltop_350_351 top350 top351 {l}
Rbot_350_351 bot350 bot351 {r}
Lbot_350_351 bot350 bot351 {l}
Rtop_350_380 top350 top380 {r}
Ltop_350_380 top350 top380 {l}
Rbot_350_380 bot350 bot380 {r}
Lbot_350_380 bot350 bot380 {l}
C350 top350 bot350 {c}
Rtop_351_352 top351 top352 {r}
Ltop_351_352 top351 top352 {l}
Rbot_351_352 bot351 bot352 {r}
Lbot_351_352 bot351 bot352 {l}
Rtop_351_381 top351 top381 {r}
Ltop_351_381 top351 top381 {l}
Rbot_351_381 bot351 bot381 {r}
Lbot_351_381 bot351 bot381 {l}
C351 top351 bot351 {c}
Rtop_352_353 top352 top353 {r}
Ltop_352_353 top352 top353 {l}
Rbot_352_353 bot352 bot353 {r}
Lbot_352_353 bot352 bot353 {l}
Rtop_352_382 top352 top382 {r}
Ltop_352_382 top352 top382 {l}
Rbot_352_382 bot352 bot382 {r}
Lbot_352_382 bot352 bot382 {l}
C352 top352 bot352 {c}
Rtop_353_354 top353 top354 {r}
Ltop_353_354 top353 top354 {l}
Rbot_353_354 bot353 bot354 {r}
Lbot_353_354 bot353 bot354 {l}
Rtop_353_383 top353 top383 {r}
Ltop_353_383 top353 top383 {l}
Rbot_353_383 bot353 bot383 {r}
Lbot_353_383 bot353 bot383 {l}
C353 top353 bot353 {c}
Rtop_354_355 top354 top355 {r}
Ltop_354_355 top354 top355 {l}
Rbot_354_355 bot354 bot355 {r}
Lbot_354_355 bot354 bot355 {l}
Rtop_354_384 top354 top384 {r}
Ltop_354_384 top354 top384 {l}
Rbot_354_384 bot354 bot384 {r}
Lbot_354_384 bot354 bot384 {l}
C354 top354 bot354 {c}
Rtop_355_356 top355 top356 {r}
Ltop_355_356 top355 top356 {l}
Rbot_355_356 bot355 bot356 {r}
Lbot_355_356 bot355 bot356 {l}
Rtop_355_385 top355 top385 {r}
Ltop_355_385 top355 top385 {l}
Rbot_355_385 bot355 bot385 {r}
Lbot_355_385 bot355 bot385 {l}
C355 top355 bot355 {c}
Rtop_356_357 top356 top357 {r}
Ltop_356_357 top356 top357 {l}
Rbot_356_357 bot356 bot357 {r}
Lbot_356_357 bot356 bot357 {l}
Rtop_356_386 top356 top386 {r}
Ltop_356_386 top356 top386 {l}
Rbot_356_386 bot356 bot386 {r}
Lbot_356_386 bot356 bot386 {l}
C356 top356 bot356 {c}
Rtop_357_358 top357 top358 {r}
Ltop_357_358 top357 top358 {l}
Rbot_357_358 bot357 bot358 {r}
Lbot_357_358 bot357 bot358 {l}
Rtop_357_387 top357 top387 {r}
Ltop_357_387 top357 top387 {l}
Rbot_357_387 bot357 bot387 {r}
Lbot_357_387 bot357 bot387 {l}
C357 top357 bot357 {c}
Rtop_358_359 top358 top359 {r}
Ltop_358_359 top358 top359 {l}
Rbot_358_359 bot358 bot359 {r}
Lbot_358_359 bot358 bot359 {l}
Rtop_358_388 top358 top388 {r}
Ltop_358_388 top358 top388 {l}
Rbot_358_388 bot358 bot388 {r}
Lbot_358_388 bot358 bot388 {l}
C358 top358 bot358 {c}
Rtop_359_360 top359 top360 {r}
Ltop_359_360 top359 top360 {l}
Rbot_359_360 bot359 bot360 {r}
Lbot_359_360 bot359 bot360 {l}
Rtop_359_389 top359 top389 {r}
Ltop_359_389 top359 top389 {l}
Rbot_359_389 bot359 bot389 {r}
Lbot_359_389 bot359 bot389 {l}
C359 top359 bot359 {c}
Rtop_360_390 top360 top390 {r}
Ltop_360_390 top360 top390 {l}
Rbot_360_390 bot360 bot390 {r}
Lbot_360_390 bot360 bot390 {l}
C360 top360 bot360 {c}
Rtop_361_362 top361 top362 {r}
Ltop_361_362 top361 top362 {l}
Rbot_361_362 bot361 bot362 {r}
Lbot_361_362 bot361 bot362 {l}
Rtop_361_391 top361 top391 {r}
Ltop_361_391 top361 top391 {l}
Rbot_361_391 bot361 bot391 {r}
Lbot_361_391 bot361 bot391 {l}
C361 top361 bot361 {c}
Rtop_362_363 top362 top363 {r}
Ltop_362_363 top362 top363 {l}
Rbot_362_363 bot362 bot363 {r}
Lbot_362_363 bot362 bot363 {l}
Rtop_362_392 top362 top392 {r}
Ltop_362_392 top362 top392 {l}
Rbot_362_392 bot362 bot392 {r}
Lbot_362_392 bot362 bot392 {l}
C362 top362 bot362 {c}
Rtop_363_364 top363 top364 {r}
Ltop_363_364 top363 top364 {l}
Rbot_363_364 bot363 bot364 {r}
Lbot_363_364 bot363 bot364 {l}
Rtop_363_393 top363 top393 {r}
Ltop_363_393 top363 top393 {l}
Rbot_363_393 bot363 bot393 {r}
Lbot_363_393 bot363 bot393 {l}
C363 top363 bot363 {c}
Rtop_364_365 top364 top365 {r}
Ltop_364_365 top364 top365 {l}
Rbot_364_365 bot364 bot365 {r}
Lbot_364_365 bot364 bot365 {l}
Rtop_364_394 top364 top394 {r}
Ltop_364_394 top364 top394 {l}
Rbot_364_394 bot364 bot394 {r}
Lbot_364_394 bot364 bot394 {l}
C364 top364 bot364 {c}
Rtop_365_366 top365 top366 {r}
Ltop_365_366 top365 top366 {l}
Rbot_365_366 bot365 bot366 {r}
Lbot_365_366 bot365 bot366 {l}
Rtop_365_395 top365 top395 {r}
Ltop_365_395 top365 top395 {l}
Rbot_365_395 bot365 bot395 {r}
Lbot_365_395 bot365 bot395 {l}
C365 top365 bot365 {c}
Rtop_366_367 top366 top367 {r}
Ltop_366_367 top366 top367 {l}
Rbot_366_367 bot366 bot367 {r}
Lbot_366_367 bot366 bot367 {l}
Rtop_366_396 top366 top396 {r}
Ltop_366_396 top366 top396 {l}
Rbot_366_396 bot366 bot396 {r}
Lbot_366_396 bot366 bot396 {l}
C366 top366 bot366 {c}
Rtop_367_368 top367 top368 {r}
Ltop_367_368 top367 top368 {l}
Rbot_367_368 bot367 bot368 {r}
Lbot_367_368 bot367 bot368 {l}
Rtop_367_397 top367 top397 {r}
Ltop_367_397 top367 top397 {l}
Rbot_367_397 bot367 bot397 {r}
Lbot_367_397 bot367 bot397 {l}
C367 top367 bot367 {c}
Rtop_368_369 top368 top369 {r}
Ltop_368_369 top368 top369 {l}
Rbot_368_369 bot368 bot369 {r}
Lbot_368_369 bot368 bot369 {l}
Rtop_368_398 top368 top398 {r}
Ltop_368_398 top368 top398 {l}
Rbot_368_398 bot368 bot398 {r}
Lbot_368_398 bot368 bot398 {l}
C368 top368 bot368 {c}
Rtop_369_370 top369 top370 {r}
Ltop_369_370 top369 top370 {l}
Rbot_369_370 bot369 bot370 {r}
Lbot_369_370 bot369 bot370 {l}
Rtop_369_399 top369 top399 {r}
Ltop_369_399 top369 top399 {l}
Rbot_369_399 bot369 bot399 {r}
Lbot_369_399 bot369 bot399 {l}
C369 top369 bot369 {c}
Rtop_370_371 top370 top371 {r}
Ltop_370_371 top370 top371 {l}
Rbot_370_371 bot370 bot371 {r}
Lbot_370_371 bot370 bot371 {l}
Rtop_370_400 top370 top400 {r}
Ltop_370_400 top370 top400 {l}
Rbot_370_400 bot370 bot400 {r}
Lbot_370_400 bot370 bot400 {l}
C370 top370 bot370 {c}
Rtop_371_372 top371 top372 {r}
Ltop_371_372 top371 top372 {l}
Rbot_371_372 bot371 bot372 {r}
Lbot_371_372 bot371 bot372 {l}
Rtop_371_401 top371 top401 {r}
Ltop_371_401 top371 top401 {l}
Rbot_371_401 bot371 bot401 {r}
Lbot_371_401 bot371 bot401 {l}
C371 top371 bot371 {c}
Rtop_372_373 top372 top373 {r}
Ltop_372_373 top372 top373 {l}
Rbot_372_373 bot372 bot373 {r}
Lbot_372_373 bot372 bot373 {l}
Rtop_372_402 top372 top402 {r}
Ltop_372_402 top372 top402 {l}
Rbot_372_402 bot372 bot402 {r}
Lbot_372_402 bot372 bot402 {l}
C372 top372 bot372 {c}
Rtop_373_374 top373 top374 {r}
Ltop_373_374 top373 top374 {l}
Rbot_373_374 bot373 bot374 {r}
Lbot_373_374 bot373 bot374 {l}
Rtop_373_403 top373 top403 {r}
Ltop_373_403 top373 top403 {l}
Rbot_373_403 bot373 bot403 {r}
Lbot_373_403 bot373 bot403 {l}
C373 top373 bot373 {c}
Rtop_374_375 top374 top375 {r}
Ltop_374_375 top374 top375 {l}
Rbot_374_375 bot374 bot375 {r}
Lbot_374_375 bot374 bot375 {l}
Rtop_374_404 top374 top404 {r}
Ltop_374_404 top374 top404 {l}
Rbot_374_404 bot374 bot404 {r}
Lbot_374_404 bot374 bot404 {l}
C374 top374 bot374 {c}
Rtop_375_376 top375 top376 {r}
Ltop_375_376 top375 top376 {l}
Rbot_375_376 bot375 bot376 {r}
Lbot_375_376 bot375 bot376 {l}
Rtop_375_405 top375 top405 {r}
Ltop_375_405 top375 top405 {l}
Rbot_375_405 bot375 bot405 {r}
Lbot_375_405 bot375 bot405 {l}
C375 top375 bot375 {c}
Rtop_376_377 top376 top377 {r}
Ltop_376_377 top376 top377 {l}
Rbot_376_377 bot376 bot377 {r}
Lbot_376_377 bot376 bot377 {l}
Rtop_376_406 top376 top406 {r}
Ltop_376_406 top376 top406 {l}
Rbot_376_406 bot376 bot406 {r}
Lbot_376_406 bot376 bot406 {l}
C376 top376 bot376 {c}
Rtop_377_378 top377 top378 {r}
Ltop_377_378 top377 top378 {l}
Rbot_377_378 bot377 bot378 {r}
Lbot_377_378 bot377 bot378 {l}
Rtop_377_407 top377 top407 {r}
Ltop_377_407 top377 top407 {l}
Rbot_377_407 bot377 bot407 {r}
Lbot_377_407 bot377 bot407 {l}
C377 top377 bot377 {c}
Rtop_378_379 top378 top379 {r}
Ltop_378_379 top378 top379 {l}
Rbot_378_379 bot378 bot379 {r}
Lbot_378_379 bot378 bot379 {l}
Rtop_378_408 top378 top408 {r}
Ltop_378_408 top378 top408 {l}
Rbot_378_408 bot378 bot408 {r}
Lbot_378_408 bot378 bot408 {l}
C378 top378 bot378 {c}
Rtop_379_380 top379 top380 {r}
Ltop_379_380 top379 top380 {l}
Rbot_379_380 bot379 bot380 {r}
Lbot_379_380 bot379 bot380 {l}
Rtop_379_409 top379 top409 {r}
Ltop_379_409 top379 top409 {l}
Rbot_379_409 bot379 bot409 {r}
Lbot_379_409 bot379 bot409 {l}
C379 top379 bot379 {c}
Rtop_380_381 top380 top381 {r}
Ltop_380_381 top380 top381 {l}
Rbot_380_381 bot380 bot381 {r}
Lbot_380_381 bot380 bot381 {l}
Rtop_380_410 top380 top410 {r}
Ltop_380_410 top380 top410 {l}
Rbot_380_410 bot380 bot410 {r}
Lbot_380_410 bot380 bot410 {l}
C380 top380 bot380 {c}
Rtop_381_382 top381 top382 {r}
Ltop_381_382 top381 top382 {l}
Rbot_381_382 bot381 bot382 {r}
Lbot_381_382 bot381 bot382 {l}
Rtop_381_411 top381 top411 {r}
Ltop_381_411 top381 top411 {l}
Rbot_381_411 bot381 bot411 {r}
Lbot_381_411 bot381 bot411 {l}
C381 top381 bot381 {c}
Rtop_382_383 top382 top383 {r}
Ltop_382_383 top382 top383 {l}
Rbot_382_383 bot382 bot383 {r}
Lbot_382_383 bot382 bot383 {l}
Rtop_382_412 top382 top412 {r}
Ltop_382_412 top382 top412 {l}
Rbot_382_412 bot382 bot412 {r}
Lbot_382_412 bot382 bot412 {l}
C382 top382 bot382 {c}
Rtop_383_384 top383 top384 {r}
Ltop_383_384 top383 top384 {l}
Rbot_383_384 bot383 bot384 {r}
Lbot_383_384 bot383 bot384 {l}
Rtop_383_413 top383 top413 {r}
Ltop_383_413 top383 top413 {l}
Rbot_383_413 bot383 bot413 {r}
Lbot_383_413 bot383 bot413 {l}
C383 top383 bot383 {c}
Rtop_384_385 top384 top385 {r}
Ltop_384_385 top384 top385 {l}
Rbot_384_385 bot384 bot385 {r}
Lbot_384_385 bot384 bot385 {l}
Rtop_384_414 top384 top414 {r}
Ltop_384_414 top384 top414 {l}
Rbot_384_414 bot384 bot414 {r}
Lbot_384_414 bot384 bot414 {l}
C384 top384 bot384 {c}
Rtop_385_386 top385 top386 {r}
Ltop_385_386 top385 top386 {l}
Rbot_385_386 bot385 bot386 {r}
Lbot_385_386 bot385 bot386 {l}
Rtop_385_415 top385 top415 {r}
Ltop_385_415 top385 top415 {l}
Rbot_385_415 bot385 bot415 {r}
Lbot_385_415 bot385 bot415 {l}
C385 top385 bot385 {c}
Rtop_386_387 top386 top387 {r}
Ltop_386_387 top386 top387 {l}
Rbot_386_387 bot386 bot387 {r}
Lbot_386_387 bot386 bot387 {l}
Rtop_386_416 top386 top416 {r}
Ltop_386_416 top386 top416 {l}
Rbot_386_416 bot386 bot416 {r}
Lbot_386_416 bot386 bot416 {l}
C386 top386 bot386 {c}
Rtop_387_388 top387 top388 {r}
Ltop_387_388 top387 top388 {l}
Rbot_387_388 bot387 bot388 {r}
Lbot_387_388 bot387 bot388 {l}
Rtop_387_417 top387 top417 {r}
Ltop_387_417 top387 top417 {l}
Rbot_387_417 bot387 bot417 {r}
Lbot_387_417 bot387 bot417 {l}
C387 top387 bot387 {c}
Rtop_388_389 top388 top389 {r}
Ltop_388_389 top388 top389 {l}
Rbot_388_389 bot388 bot389 {r}
Lbot_388_389 bot388 bot389 {l}
Rtop_388_418 top388 top418 {r}
Ltop_388_418 top388 top418 {l}
Rbot_388_418 bot388 bot418 {r}
Lbot_388_418 bot388 bot418 {l}
C388 top388 bot388 {c}
Rtop_389_390 top389 top390 {r}
Ltop_389_390 top389 top390 {l}
Rbot_389_390 bot389 bot390 {r}
Lbot_389_390 bot389 bot390 {l}
Rtop_389_419 top389 top419 {r}
Ltop_389_419 top389 top419 {l}
Rbot_389_419 bot389 bot419 {r}
Lbot_389_419 bot389 bot419 {l}
C389 top389 bot389 {c}
Rtop_390_420 top390 top420 {r}
Ltop_390_420 top390 top420 {l}
Rbot_390_420 bot390 bot420 {r}
Lbot_390_420 bot390 bot420 {l}
C390 top390 bot390 {c}
Rtop_391_392 top391 top392 {r}
Ltop_391_392 top391 top392 {l}
Rbot_391_392 bot391 bot392 {r}
Lbot_391_392 bot391 bot392 {l}
Rtop_391_421 top391 top421 {r}
Ltop_391_421 top391 top421 {l}
Rbot_391_421 bot391 bot421 {r}
Lbot_391_421 bot391 bot421 {l}
C391 top391 bot391 {c}
Rtop_392_393 top392 top393 {r}
Ltop_392_393 top392 top393 {l}
Rbot_392_393 bot392 bot393 {r}
Lbot_392_393 bot392 bot393 {l}
Rtop_392_422 top392 top422 {r}
Ltop_392_422 top392 top422 {l}
Rbot_392_422 bot392 bot422 {r}
Lbot_392_422 bot392 bot422 {l}
C392 top392 bot392 {c}
Rtop_393_394 top393 top394 {r}
Ltop_393_394 top393 top394 {l}
Rbot_393_394 bot393 bot394 {r}
Lbot_393_394 bot393 bot394 {l}
Rtop_393_423 top393 top423 {r}
Ltop_393_423 top393 top423 {l}
Rbot_393_423 bot393 bot423 {r}
Lbot_393_423 bot393 bot423 {l}
C393 top393 bot393 {c}
Rtop_394_395 top394 top395 {r}
Ltop_394_395 top394 top395 {l}
Rbot_394_395 bot394 bot395 {r}
Lbot_394_395 bot394 bot395 {l}
Rtop_394_424 top394 top424 {r}
Ltop_394_424 top394 top424 {l}
Rbot_394_424 bot394 bot424 {r}
Lbot_394_424 bot394 bot424 {l}
C394 top394 bot394 {c}
Rtop_395_396 top395 top396 {r}
Ltop_395_396 top395 top396 {l}
Rbot_395_396 bot395 bot396 {r}
Lbot_395_396 bot395 bot396 {l}
Rtop_395_425 top395 top425 {r}
Ltop_395_425 top395 top425 {l}
Rbot_395_425 bot395 bot425 {r}
Lbot_395_425 bot395 bot425 {l}
C395 top395 bot395 {c}
Rtop_396_397 top396 top397 {r}
Ltop_396_397 top396 top397 {l}
Rbot_396_397 bot396 bot397 {r}
Lbot_396_397 bot396 bot397 {l}
Rtop_396_426 top396 top426 {r}
Ltop_396_426 top396 top426 {l}
Rbot_396_426 bot396 bot426 {r}
Lbot_396_426 bot396 bot426 {l}
C396 top396 bot396 {c}
Rtop_397_398 top397 top398 {r}
Ltop_397_398 top397 top398 {l}
Rbot_397_398 bot397 bot398 {r}
Lbot_397_398 bot397 bot398 {l}
Rtop_397_427 top397 top427 {r}
Ltop_397_427 top397 top427 {l}
Rbot_397_427 bot397 bot427 {r}
Lbot_397_427 bot397 bot427 {l}
C397 top397 bot397 {c}
Rtop_398_399 top398 top399 {r}
Ltop_398_399 top398 top399 {l}
Rbot_398_399 bot398 bot399 {r}
Lbot_398_399 bot398 bot399 {l}
Rtop_398_428 top398 top428 {r}
Ltop_398_428 top398 top428 {l}
Rbot_398_428 bot398 bot428 {r}
Lbot_398_428 bot398 bot428 {l}
C398 top398 bot398 {c}
Rtop_399_400 top399 top400 {r}
Ltop_399_400 top399 top400 {l}
Rbot_399_400 bot399 bot400 {r}
Lbot_399_400 bot399 bot400 {l}
Rtop_399_429 top399 top429 {r}
Ltop_399_429 top399 top429 {l}
Rbot_399_429 bot399 bot429 {r}
Lbot_399_429 bot399 bot429 {l}
C399 top399 bot399 {c}
Rtop_400_401 top400 top401 {r}
Ltop_400_401 top400 top401 {l}
Rbot_400_401 bot400 bot401 {r}
Lbot_400_401 bot400 bot401 {l}
Rtop_400_430 top400 top430 {r}
Ltop_400_430 top400 top430 {l}
Rbot_400_430 bot400 bot430 {r}
Lbot_400_430 bot400 bot430 {l}
C400 top400 bot400 {c}
Rtop_401_402 top401 top402 {r}
Ltop_401_402 top401 top402 {l}
Rbot_401_402 bot401 bot402 {r}
Lbot_401_402 bot401 bot402 {l}
Rtop_401_431 top401 top431 {r}
Ltop_401_431 top401 top431 {l}
Rbot_401_431 bot401 bot431 {r}
Lbot_401_431 bot401 bot431 {l}
C401 top401 bot401 {c}
Rtop_402_403 top402 top403 {r}
Ltop_402_403 top402 top403 {l}
Rbot_402_403 bot402 bot403 {r}
Lbot_402_403 bot402 bot403 {l}
Rtop_402_432 top402 top432 {r}
Ltop_402_432 top402 top432 {l}
Rbot_402_432 bot402 bot432 {r}
Lbot_402_432 bot402 bot432 {l}
C402 top402 bot402 {c}
Rtop_403_404 top403 top404 {r}
Ltop_403_404 top403 top404 {l}
Rbot_403_404 bot403 bot404 {r}
Lbot_403_404 bot403 bot404 {l}
Rtop_403_433 top403 top433 {r}
Ltop_403_433 top403 top433 {l}
Rbot_403_433 bot403 bot433 {r}
Lbot_403_433 bot403 bot433 {l}
C403 top403 bot403 {c}
Rtop_404_405 top404 top405 {r}
Ltop_404_405 top404 top405 {l}
Rbot_404_405 bot404 bot405 {r}
Lbot_404_405 bot404 bot405 {l}
Rtop_404_434 top404 top434 {r}
Ltop_404_434 top404 top434 {l}
Rbot_404_434 bot404 bot434 {r}
Lbot_404_434 bot404 bot434 {l}
C404 top404 bot404 {c}
Rtop_405_406 top405 top406 {r}
Ltop_405_406 top405 top406 {l}
Rbot_405_406 bot405 bot406 {r}
Lbot_405_406 bot405 bot406 {l}
Rtop_405_435 top405 top435 {r}
Ltop_405_435 top405 top435 {l}
Rbot_405_435 bot405 bot435 {r}
Lbot_405_435 bot405 bot435 {l}
C405 top405 bot405 {c}
Rtop_406_407 top406 top407 {r}
Ltop_406_407 top406 top407 {l}
Rbot_406_407 bot406 bot407 {r}
Lbot_406_407 bot406 bot407 {l}
Rtop_406_436 top406 top436 {r}
Ltop_406_436 top406 top436 {l}
Rbot_406_436 bot406 bot436 {r}
Lbot_406_436 bot406 bot436 {l}
C406 top406 bot406 {c}
Rtop_407_408 top407 top408 {r}
Ltop_407_408 top407 top408 {l}
Rbot_407_408 bot407 bot408 {r}
Lbot_407_408 bot407 bot408 {l}
Rtop_407_437 top407 top437 {r}
Ltop_407_437 top407 top437 {l}
Rbot_407_437 bot407 bot437 {r}
Lbot_407_437 bot407 bot437 {l}
C407 top407 bot407 {c}
Rtop_408_409 top408 top409 {r}
Ltop_408_409 top408 top409 {l}
Rbot_408_409 bot408 bot409 {r}
Lbot_408_409 bot408 bot409 {l}
Rtop_408_438 top408 top438 {r}
Ltop_408_438 top408 top438 {l}
Rbot_408_438 bot408 bot438 {r}
Lbot_408_438 bot408 bot438 {l}
C408 top408 bot408 {c}
Rtop_409_410 top409 top410 {r}
Ltop_409_410 top409 top410 {l}
Rbot_409_410 bot409 bot410 {r}
Lbot_409_410 bot409 bot410 {l}
Rtop_409_439 top409 top439 {r}
Ltop_409_439 top409 top439 {l}
Rbot_409_439 bot409 bot439 {r}
Lbot_409_439 bot409 bot439 {l}
C409 top409 bot409 {c}
Rtop_410_411 top410 top411 {r}
Ltop_410_411 top410 top411 {l}
Rbot_410_411 bot410 bot411 {r}
Lbot_410_411 bot410 bot411 {l}
Rtop_410_440 top410 top440 {r}
Ltop_410_440 top410 top440 {l}
Rbot_410_440 bot410 bot440 {r}
Lbot_410_440 bot410 bot440 {l}
C410 top410 bot410 {c}
Rtop_411_412 top411 top412 {r}
Ltop_411_412 top411 top412 {l}
Rbot_411_412 bot411 bot412 {r}
Lbot_411_412 bot411 bot412 {l}
Rtop_411_441 top411 top441 {r}
Ltop_411_441 top411 top441 {l}
Rbot_411_441 bot411 bot441 {r}
Lbot_411_441 bot411 bot441 {l}
C411 top411 bot411 {c}
Rtop_412_413 top412 top413 {r}
Ltop_412_413 top412 top413 {l}
Rbot_412_413 bot412 bot413 {r}
Lbot_412_413 bot412 bot413 {l}
Rtop_412_442 top412 top442 {r}
Ltop_412_442 top412 top442 {l}
Rbot_412_442 bot412 bot442 {r}
Lbot_412_442 bot412 bot442 {l}
C412 top412 bot412 {c}
Rtop_413_414 top413 top414 {r}
Ltop_413_414 top413 top414 {l}
Rbot_413_414 bot413 bot414 {r}
Lbot_413_414 bot413 bot414 {l}
Rtop_413_443 top413 top443 {r}
Ltop_413_443 top413 top443 {l}
Rbot_413_443 bot413 bot443 {r}
Lbot_413_443 bot413 bot443 {l}
C413 top413 bot413 {c}
Rtop_414_415 top414 top415 {r}
Ltop_414_415 top414 top415 {l}
Rbot_414_415 bot414 bot415 {r}
Lbot_414_415 bot414 bot415 {l}
Rtop_414_444 top414 top444 {r}
Ltop_414_444 top414 top444 {l}
Rbot_414_444 bot414 bot444 {r}
Lbot_414_444 bot414 bot444 {l}
C414 top414 bot414 {c}
Rtop_415_416 top415 top416 {r}
Ltop_415_416 top415 top416 {l}
Rbot_415_416 bot415 bot416 {r}
Lbot_415_416 bot415 bot416 {l}
Rtop_415_445 top415 top445 {r}
Ltop_415_445 top415 top445 {l}
Rbot_415_445 bot415 bot445 {r}
Lbot_415_445 bot415 bot445 {l}
C415 top415 bot415 {c}
Rtop_416_417 top416 top417 {r}
Ltop_416_417 top416 top417 {l}
Rbot_416_417 bot416 bot417 {r}
Lbot_416_417 bot416 bot417 {l}
Rtop_416_446 top416 top446 {r}
Ltop_416_446 top416 top446 {l}
Rbot_416_446 bot416 bot446 {r}
Lbot_416_446 bot416 bot446 {l}
C416 top416 bot416 {c}
Rtop_417_418 top417 top418 {r}
Ltop_417_418 top417 top418 {l}
Rbot_417_418 bot417 bot418 {r}
Lbot_417_418 bot417 bot418 {l}
Rtop_417_447 top417 top447 {r}
Ltop_417_447 top417 top447 {l}
Rbot_417_447 bot417 bot447 {r}
Lbot_417_447 bot417 bot447 {l}
C417 top417 bot417 {c}
Rtop_418_419 top418 top419 {r}
Ltop_418_419 top418 top419 {l}
Rbot_418_419 bot418 bot419 {r}
Lbot_418_419 bot418 bot419 {l}
Rtop_418_448 top418 top448 {r}
Ltop_418_448 top418 top448 {l}
Rbot_418_448 bot418 bot448 {r}
Lbot_418_448 bot418 bot448 {l}
C418 top418 bot418 {c}
Rtop_419_420 top419 top420 {r}
Ltop_419_420 top419 top420 {l}
Rbot_419_420 bot419 bot420 {r}
Lbot_419_420 bot419 bot420 {l}
Rtop_419_449 top419 top449 {r}
Ltop_419_449 top419 top449 {l}
Rbot_419_449 bot419 bot449 {r}
Lbot_419_449 bot419 bot449 {l}
C419 top419 bot419 {c}
Rtop_420_450 top420 top450 {r}
Ltop_420_450 top420 top450 {l}
Rbot_420_450 bot420 bot450 {r}
Lbot_420_450 bot420 bot450 {l}
C420 top420 bot420 {c}
Rtop_421_422 top421 top422 {r}
Ltop_421_422 top421 top422 {l}
Rbot_421_422 bot421 bot422 {r}
Lbot_421_422 bot421 bot422 {l}
Rtop_421_451 top421 top451 {r}
Ltop_421_451 top421 top451 {l}
Rbot_421_451 bot421 bot451 {r}
Lbot_421_451 bot421 bot451 {l}
C421 top421 bot421 {c}
Rtop_422_423 top422 top423 {r}
Ltop_422_423 top422 top423 {l}
Rbot_422_423 bot422 bot423 {r}
Lbot_422_423 bot422 bot423 {l}
Rtop_422_452 top422 top452 {r}
Ltop_422_452 top422 top452 {l}
Rbot_422_452 bot422 bot452 {r}
Lbot_422_452 bot422 bot452 {l}
C422 top422 bot422 {c}
Rtop_423_424 top423 top424 {r}
Ltop_423_424 top423 top424 {l}
Rbot_423_424 bot423 bot424 {r}
Lbot_423_424 bot423 bot424 {l}
Rtop_423_453 top423 top453 {r}
Ltop_423_453 top423 top453 {l}
Rbot_423_453 bot423 bot453 {r}
Lbot_423_453 bot423 bot453 {l}
C423 top423 bot423 {c}
Rtop_424_425 top424 top425 {r}
Ltop_424_425 top424 top425 {l}
Rbot_424_425 bot424 bot425 {r}
Lbot_424_425 bot424 bot425 {l}
Rtop_424_454 top424 top454 {r}
Ltop_424_454 top424 top454 {l}
Rbot_424_454 bot424 bot454 {r}
Lbot_424_454 bot424 bot454 {l}
C424 top424 bot424 {c}
Rtop_425_426 top425 top426 {r}
Ltop_425_426 top425 top426 {l}
Rbot_425_426 bot425 bot426 {r}
Lbot_425_426 bot425 bot426 {l}
Rtop_425_455 top425 top455 {r}
Ltop_425_455 top425 top455 {l}
Rbot_425_455 bot425 bot455 {r}
Lbot_425_455 bot425 bot455 {l}
C425 top425 bot425 {c}
Rtop_426_427 top426 top427 {r}
Ltop_426_427 top426 top427 {l}
Rbot_426_427 bot426 bot427 {r}
Lbot_426_427 bot426 bot427 {l}
Rtop_426_456 top426 top456 {r}
Ltop_426_456 top426 top456 {l}
Rbot_426_456 bot426 bot456 {r}
Lbot_426_456 bot426 bot456 {l}
C426 top426 bot426 {c}
Rtop_427_428 top427 top428 {r}
Ltop_427_428 top427 top428 {l}
Rbot_427_428 bot427 bot428 {r}
Lbot_427_428 bot427 bot428 {l}
Rtop_427_457 top427 top457 {r}
Ltop_427_457 top427 top457 {l}
Rbot_427_457 bot427 bot457 {r}
Lbot_427_457 bot427 bot457 {l}
C427 top427 bot427 {c}
Rtop_428_429 top428 top429 {r}
Ltop_428_429 top428 top429 {l}
Rbot_428_429 bot428 bot429 {r}
Lbot_428_429 bot428 bot429 {l}
Rtop_428_458 top428 top458 {r}
Ltop_428_458 top428 top458 {l}
Rbot_428_458 bot428 bot458 {r}
Lbot_428_458 bot428 bot458 {l}
C428 top428 bot428 {c}
Rtop_429_430 top429 top430 {r}
Ltop_429_430 top429 top430 {l}
Rbot_429_430 bot429 bot430 {r}
Lbot_429_430 bot429 bot430 {l}
Rtop_429_459 top429 top459 {r}
Ltop_429_459 top429 top459 {l}
Rbot_429_459 bot429 bot459 {r}
Lbot_429_459 bot429 bot459 {l}
C429 top429 bot429 {c}
Rtop_430_431 top430 top431 {r}
Ltop_430_431 top430 top431 {l}
Rbot_430_431 bot430 bot431 {r}
Lbot_430_431 bot430 bot431 {l}
Rtop_430_460 top430 top460 {r}
Ltop_430_460 top430 top460 {l}
Rbot_430_460 bot430 bot460 {r}
Lbot_430_460 bot430 bot460 {l}
C430 top430 bot430 {c}
Rtop_431_432 top431 top432 {r}
Ltop_431_432 top431 top432 {l}
Rbot_431_432 bot431 bot432 {r}
Lbot_431_432 bot431 bot432 {l}
Rtop_431_461 top431 top461 {r}
Ltop_431_461 top431 top461 {l}
Rbot_431_461 bot431 bot461 {r}
Lbot_431_461 bot431 bot461 {l}
C431 top431 bot431 {c}
Rtop_432_433 top432 top433 {r}
Ltop_432_433 top432 top433 {l}
Rbot_432_433 bot432 bot433 {r}
Lbot_432_433 bot432 bot433 {l}
Rtop_432_462 top432 top462 {r}
Ltop_432_462 top432 top462 {l}
Rbot_432_462 bot432 bot462 {r}
Lbot_432_462 bot432 bot462 {l}
C432 top432 bot432 {c}
Rtop_433_434 top433 top434 {r}
Ltop_433_434 top433 top434 {l}
Rbot_433_434 bot433 bot434 {r}
Lbot_433_434 bot433 bot434 {l}
Rtop_433_463 top433 top463 {r}
Ltop_433_463 top433 top463 {l}
Rbot_433_463 bot433 bot463 {r}
Lbot_433_463 bot433 bot463 {l}
C433 top433 bot433 {c}
Rtop_434_435 top434 top435 {r}
Ltop_434_435 top434 top435 {l}
Rbot_434_435 bot434 bot435 {r}
Lbot_434_435 bot434 bot435 {l}
Rtop_434_464 top434 top464 {r}
Ltop_434_464 top434 top464 {l}
Rbot_434_464 bot434 bot464 {r}
Lbot_434_464 bot434 bot464 {l}
C434 top434 bot434 {c}
Rtop_435_436 top435 top436 {r}
Ltop_435_436 top435 top436 {l}
Rbot_435_436 bot435 bot436 {r}
Lbot_435_436 bot435 bot436 {l}
Rtop_435_465 top435 top465 {r}
Ltop_435_465 top435 top465 {l}
Rbot_435_465 bot435 bot465 {r}
Lbot_435_465 bot435 bot465 {l}
C435 top435 bot435 {c}
Rtop_436_437 top436 top437 {r}
Ltop_436_437 top436 top437 {l}
Rbot_436_437 bot436 bot437 {r}
Lbot_436_437 bot436 bot437 {l}
Rtop_436_466 top436 top466 {r}
Ltop_436_466 top436 top466 {l}
Rbot_436_466 bot436 bot466 {r}
Lbot_436_466 bot436 bot466 {l}
C436 top436 bot436 {c}
Rtop_437_438 top437 top438 {r}
Ltop_437_438 top437 top438 {l}
Rbot_437_438 bot437 bot438 {r}
Lbot_437_438 bot437 bot438 {l}
Rtop_437_467 top437 top467 {r}
Ltop_437_467 top437 top467 {l}
Rbot_437_467 bot437 bot467 {r}
Lbot_437_467 bot437 bot467 {l}
C437 top437 bot437 {c}
Rtop_438_439 top438 top439 {r}
Ltop_438_439 top438 top439 {l}
Rbot_438_439 bot438 bot439 {r}
Lbot_438_439 bot438 bot439 {l}
Rtop_438_468 top438 top468 {r}
Ltop_438_468 top438 top468 {l}
Rbot_438_468 bot438 bot468 {r}
Lbot_438_468 bot438 bot468 {l}
C438 top438 bot438 {c}
Rtop_439_440 top439 top440 {r}
Ltop_439_440 top439 top440 {l}
Rbot_439_440 bot439 bot440 {r}
Lbot_439_440 bot439 bot440 {l}
Rtop_439_469 top439 top469 {r}
Ltop_439_469 top439 top469 {l}
Rbot_439_469 bot439 bot469 {r}
Lbot_439_469 bot439 bot469 {l}
C439 top439 bot439 {c}
Rtop_440_441 top440 top441 {r}
Ltop_440_441 top440 top441 {l}
Rbot_440_441 bot440 bot441 {r}
Lbot_440_441 bot440 bot441 {l}
Rtop_440_470 top440 top470 {r}
Ltop_440_470 top440 top470 {l}
Rbot_440_470 bot440 bot470 {r}
Lbot_440_470 bot440 bot470 {l}
C440 top440 bot440 {c}
Rtop_441_442 top441 top442 {r}
Ltop_441_442 top441 top442 {l}
Rbot_441_442 bot441 bot442 {r}
Lbot_441_442 bot441 bot442 {l}
Rtop_441_471 top441 top471 {r}
Ltop_441_471 top441 top471 {l}
Rbot_441_471 bot441 bot471 {r}
Lbot_441_471 bot441 bot471 {l}
C441 top441 bot441 {c}
Rtop_442_443 top442 top443 {r}
Ltop_442_443 top442 top443 {l}
Rbot_442_443 bot442 bot443 {r}
Lbot_442_443 bot442 bot443 {l}
Rtop_442_472 top442 top472 {r}
Ltop_442_472 top442 top472 {l}
Rbot_442_472 bot442 bot472 {r}
Lbot_442_472 bot442 bot472 {l}
C442 top442 bot442 {c}
Rtop_443_444 top443 top444 {r}
Ltop_443_444 top443 top444 {l}
Rbot_443_444 bot443 bot444 {r}
Lbot_443_444 bot443 bot444 {l}
Rtop_443_473 top443 top473 {r}
Ltop_443_473 top443 top473 {l}
Rbot_443_473 bot443 bot473 {r}
Lbot_443_473 bot443 bot473 {l}
C443 top443 bot443 {c}
Rtop_444_445 top444 top445 {r}
Ltop_444_445 top444 top445 {l}
Rbot_444_445 bot444 bot445 {r}
Lbot_444_445 bot444 bot445 {l}
Rtop_444_474 top444 top474 {r}
Ltop_444_474 top444 top474 {l}
Rbot_444_474 bot444 bot474 {r}
Lbot_444_474 bot444 bot474 {l}
C444 top444 bot444 {c}
Rtop_445_446 top445 top446 {r}
Ltop_445_446 top445 top446 {l}
Rbot_445_446 bot445 bot446 {r}
Lbot_445_446 bot445 bot446 {l}
Rtop_445_475 top445 top475 {r}
Ltop_445_475 top445 top475 {l}
Rbot_445_475 bot445 bot475 {r}
Lbot_445_475 bot445 bot475 {l}
C445 top445 bot445 {c}
Rtop_446_447 top446 top447 {r}
Ltop_446_447 top446 top447 {l}
Rbot_446_447 bot446 bot447 {r}
Lbot_446_447 bot446 bot447 {l}
Rtop_446_476 top446 top476 {r}
Ltop_446_476 top446 top476 {l}
Rbot_446_476 bot446 bot476 {r}
Lbot_446_476 bot446 bot476 {l}
C446 top446 bot446 {c}
Rtop_447_448 top447 top448 {r}
Ltop_447_448 top447 top448 {l}
Rbot_447_448 bot447 bot448 {r}
Lbot_447_448 bot447 bot448 {l}
Rtop_447_477 top447 top477 {r}
Ltop_447_477 top447 top477 {l}
Rbot_447_477 bot447 bot477 {r}
Lbot_447_477 bot447 bot477 {l}
C447 top447 bot447 {c}
Rtop_448_449 top448 top449 {r}
Ltop_448_449 top448 top449 {l}
Rbot_448_449 bot448 bot449 {r}
Lbot_448_449 bot448 bot449 {l}
Rtop_448_478 top448 top478 {r}
Ltop_448_478 top448 top478 {l}
Rbot_448_478 bot448 bot478 {r}
Lbot_448_478 bot448 bot478 {l}
C448 top448 bot448 {c}
Rtop_449_450 top449 top450 {r}
Ltop_449_450 top449 top450 {l}
Rbot_449_450 bot449 bot450 {r}
Lbot_449_450 bot449 bot450 {l}
Rtop_449_479 top449 top479 {r}
Ltop_449_479 top449 top479 {l}
Rbot_449_479 bot449 bot479 {r}
Lbot_449_479 bot449 bot479 {l}
C449 top449 bot449 {c}
Rtop_450_480 top450 top480 {r}
Ltop_450_480 top450 top480 {l}
Rbot_450_480 bot450 bot480 {r}
Lbot_450_480 bot450 bot480 {l}
C450 top450 bot450 {c}
Rtop_451_452 top451 top452 {r}
Ltop_451_452 top451 top452 {l}
Rbot_451_452 bot451 bot452 {r}
Lbot_451_452 bot451 bot452 {l}
Rtop_451_481 top451 top481 {r}
Ltop_451_481 top451 top481 {l}
Rbot_451_481 bot451 bot481 {r}
Lbot_451_481 bot451 bot481 {l}
C451 top451 bot451 {c}
Rtop_452_453 top452 top453 {r}
Ltop_452_453 top452 top453 {l}
Rbot_452_453 bot452 bot453 {r}
Lbot_452_453 bot452 bot453 {l}
Rtop_452_482 top452 top482 {r}
Ltop_452_482 top452 top482 {l}
Rbot_452_482 bot452 bot482 {r}
Lbot_452_482 bot452 bot482 {l}
C452 top452 bot452 {c}
Rtop_453_454 top453 top454 {r}
Ltop_453_454 top453 top454 {l}
Rbot_453_454 bot453 bot454 {r}
Lbot_453_454 bot453 bot454 {l}
Rtop_453_483 top453 top483 {r}
Ltop_453_483 top453 top483 {l}
Rbot_453_483 bot453 bot483 {r}
Lbot_453_483 bot453 bot483 {l}
C453 top453 bot453 {c}
Rtop_454_455 top454 top455 {r}
Ltop_454_455 top454 top455 {l}
Rbot_454_455 bot454 bot455 {r}
Lbot_454_455 bot454 bot455 {l}
Rtop_454_484 top454 top484 {r}
Ltop_454_484 top454 top484 {l}
Rbot_454_484 bot454 bot484 {r}
Lbot_454_484 bot454 bot484 {l}
C454 top454 bot454 {c}
Rtop_455_456 top455 top456 {r}
Ltop_455_456 top455 top456 {l}
Rbot_455_456 bot455 bot456 {r}
Lbot_455_456 bot455 bot456 {l}
Rtop_455_485 top455 top485 {r}
Ltop_455_485 top455 top485 {l}
Rbot_455_485 bot455 bot485 {r}
Lbot_455_485 bot455 bot485 {l}
C455 top455 bot455 {c}
Rtop_456_457 top456 top457 {r}
Ltop_456_457 top456 top457 {l}
Rbot_456_457 bot456 bot457 {r}
Lbot_456_457 bot456 bot457 {l}
Rtop_456_486 top456 top486 {r}
Ltop_456_486 top456 top486 {l}
Rbot_456_486 bot456 bot486 {r}
Lbot_456_486 bot456 bot486 {l}
C456 top456 bot456 {c}
Rtop_457_458 top457 top458 {r}
Ltop_457_458 top457 top458 {l}
Rbot_457_458 bot457 bot458 {r}
Lbot_457_458 bot457 bot458 {l}
Rtop_457_487 top457 top487 {r}
Ltop_457_487 top457 top487 {l}
Rbot_457_487 bot457 bot487 {r}
Lbot_457_487 bot457 bot487 {l}
C457 top457 bot457 {c}
Rtop_458_459 top458 top459 {r}
Ltop_458_459 top458 top459 {l}
Rbot_458_459 bot458 bot459 {r}
Lbot_458_459 bot458 bot459 {l}
Rtop_458_488 top458 top488 {r}
Ltop_458_488 top458 top488 {l}
Rbot_458_488 bot458 bot488 {r}
Lbot_458_488 bot458 bot488 {l}
C458 top458 bot458 {c}
Rtop_459_460 top459 top460 {r}
Ltop_459_460 top459 top460 {l}
Rbot_459_460 bot459 bot460 {r}
Lbot_459_460 bot459 bot460 {l}
Rtop_459_489 top459 top489 {r}
Ltop_459_489 top459 top489 {l}
Rbot_459_489 bot459 bot489 {r}
Lbot_459_489 bot459 bot489 {l}
C459 top459 bot459 {c}
Rtop_460_461 top460 top461 {r}
Ltop_460_461 top460 top461 {l}
Rbot_460_461 bot460 bot461 {r}
Lbot_460_461 bot460 bot461 {l}
Rtop_460_490 top460 top490 {r}
Ltop_460_490 top460 top490 {l}
Rbot_460_490 bot460 bot490 {r}
Lbot_460_490 bot460 bot490 {l}
C460 top460 bot460 {c}
Rtop_461_462 top461 top462 {r}
Ltop_461_462 top461 top462 {l}
Rbot_461_462 bot461 bot462 {r}
Lbot_461_462 bot461 bot462 {l}
Rtop_461_491 top461 top491 {r}
Ltop_461_491 top461 top491 {l}
Rbot_461_491 bot461 bot491 {r}
Lbot_461_491 bot461 bot491 {l}
C461 top461 bot461 {c}
Rtop_462_463 top462 top463 {r}
Ltop_462_463 top462 top463 {l}
Rbot_462_463 bot462 bot463 {r}
Lbot_462_463 bot462 bot463 {l}
Rtop_462_492 top462 top492 {r}
Ltop_462_492 top462 top492 {l}
Rbot_462_492 bot462 bot492 {r}
Lbot_462_492 bot462 bot492 {l}
C462 top462 bot462 {c}
Rtop_463_464 top463 top464 {r}
Ltop_463_464 top463 top464 {l}
Rbot_463_464 bot463 bot464 {r}
Lbot_463_464 bot463 bot464 {l}
Rtop_463_493 top463 top493 {r}
Ltop_463_493 top463 top493 {l}
Rbot_463_493 bot463 bot493 {r}
Lbot_463_493 bot463 bot493 {l}
C463 top463 bot463 {c}
Rtop_464_465 top464 top465 {r}
Ltop_464_465 top464 top465 {l}
Rbot_464_465 bot464 bot465 {r}
Lbot_464_465 bot464 bot465 {l}
Rtop_464_494 top464 top494 {r}
Ltop_464_494 top464 top494 {l}
Rbot_464_494 bot464 bot494 {r}
Lbot_464_494 bot464 bot494 {l}
C464 top464 bot464 {c}
Rtop_465_466 top465 top466 {r}
Ltop_465_466 top465 top466 {l}
Rbot_465_466 bot465 bot466 {r}
Lbot_465_466 bot465 bot466 {l}
Rtop_465_495 top465 top495 {r}
Ltop_465_495 top465 top495 {l}
Rbot_465_495 bot465 bot495 {r}
Lbot_465_495 bot465 bot495 {l}
C465 top465 bot465 {c}
Rtop_466_467 top466 top467 {r}
Ltop_466_467 top466 top467 {l}
Rbot_466_467 bot466 bot467 {r}
Lbot_466_467 bot466 bot467 {l}
Rtop_466_496 top466 top496 {r}
Ltop_466_496 top466 top496 {l}
Rbot_466_496 bot466 bot496 {r}
Lbot_466_496 bot466 bot496 {l}
C466 top466 bot466 {c}
Rtop_467_468 top467 top468 {r}
Ltop_467_468 top467 top468 {l}
Rbot_467_468 bot467 bot468 {r}
Lbot_467_468 bot467 bot468 {l}
Rtop_467_497 top467 top497 {r}
Ltop_467_497 top467 top497 {l}
Rbot_467_497 bot467 bot497 {r}
Lbot_467_497 bot467 bot497 {l}
C467 top467 bot467 {c}
Rtop_468_469 top468 top469 {r}
Ltop_468_469 top468 top469 {l}
Rbot_468_469 bot468 bot469 {r}
Lbot_468_469 bot468 bot469 {l}
Rtop_468_498 top468 top498 {r}
Ltop_468_498 top468 top498 {l}
Rbot_468_498 bot468 bot498 {r}
Lbot_468_498 bot468 bot498 {l}
C468 top468 bot468 {c}
Rtop_469_470 top469 top470 {r}
Ltop_469_470 top469 top470 {l}
Rbot_469_470 bot469 bot470 {r}
Lbot_469_470 bot469 bot470 {l}
Rtop_469_499 top469 top499 {r}
Ltop_469_499 top469 top499 {l}
Rbot_469_499 bot469 bot499 {r}
Lbot_469_499 bot469 bot499 {l}
C469 top469 bot469 {c}
Rtop_470_471 top470 top471 {r}
Ltop_470_471 top470 top471 {l}
Rbot_470_471 bot470 bot471 {r}
Lbot_470_471 bot470 bot471 {l}
Rtop_470_500 top470 top500 {r}
Ltop_470_500 top470 top500 {l}
Rbot_470_500 bot470 bot500 {r}
Lbot_470_500 bot470 bot500 {l}
C470 top470 bot470 {c}
Rtop_471_472 top471 top472 {r}
Ltop_471_472 top471 top472 {l}
Rbot_471_472 bot471 bot472 {r}
Lbot_471_472 bot471 bot472 {l}
Rtop_471_501 top471 top501 {r}
Ltop_471_501 top471 top501 {l}
Rbot_471_501 bot471 bot501 {r}
Lbot_471_501 bot471 bot501 {l}
C471 top471 bot471 {c}
Rtop_472_473 top472 top473 {r}
Ltop_472_473 top472 top473 {l}
Rbot_472_473 bot472 bot473 {r}
Lbot_472_473 bot472 bot473 {l}
Rtop_472_502 top472 top502 {r}
Ltop_472_502 top472 top502 {l}
Rbot_472_502 bot472 bot502 {r}
Lbot_472_502 bot472 bot502 {l}
C472 top472 bot472 {c}
Rtop_473_474 top473 top474 {r}
Ltop_473_474 top473 top474 {l}
Rbot_473_474 bot473 bot474 {r}
Lbot_473_474 bot473 bot474 {l}
Rtop_473_503 top473 top503 {r}
Ltop_473_503 top473 top503 {l}
Rbot_473_503 bot473 bot503 {r}
Lbot_473_503 bot473 bot503 {l}
C473 top473 bot473 {c}
Rtop_474_475 top474 top475 {r}
Ltop_474_475 top474 top475 {l}
Rbot_474_475 bot474 bot475 {r}
Lbot_474_475 bot474 bot475 {l}
Rtop_474_504 top474 top504 {r}
Ltop_474_504 top474 top504 {l}
Rbot_474_504 bot474 bot504 {r}
Lbot_474_504 bot474 bot504 {l}
C474 top474 bot474 {c}
Rtop_475_476 top475 top476 {r}
Ltop_475_476 top475 top476 {l}
Rbot_475_476 bot475 bot476 {r}
Lbot_475_476 bot475 bot476 {l}
Rtop_475_505 top475 top505 {r}
Ltop_475_505 top475 top505 {l}
Rbot_475_505 bot475 bot505 {r}
Lbot_475_505 bot475 bot505 {l}
C475 top475 bot475 {c}
Rtop_476_477 top476 top477 {r}
Ltop_476_477 top476 top477 {l}
Rbot_476_477 bot476 bot477 {r}
Lbot_476_477 bot476 bot477 {l}
Rtop_476_506 top476 top506 {r}
Ltop_476_506 top476 top506 {l}
Rbot_476_506 bot476 bot506 {r}
Lbot_476_506 bot476 bot506 {l}
C476 top476 bot476 {c}
Rtop_477_478 top477 top478 {r}
Ltop_477_478 top477 top478 {l}
Rbot_477_478 bot477 bot478 {r}
Lbot_477_478 bot477 bot478 {l}
Rtop_477_507 top477 top507 {r}
Ltop_477_507 top477 top507 {l}
Rbot_477_507 bot477 bot507 {r}
Lbot_477_507 bot477 bot507 {l}
C477 top477 bot477 {c}
Rtop_478_479 top478 top479 {r}
Ltop_478_479 top478 top479 {l}
Rbot_478_479 bot478 bot479 {r}
Lbot_478_479 bot478 bot479 {l}
Rtop_478_508 top478 top508 {r}
Ltop_478_508 top478 top508 {l}
Rbot_478_508 bot478 bot508 {r}
Lbot_478_508 bot478 bot508 {l}
C478 top478 bot478 {c}
Rtop_479_480 top479 top480 {r}
Ltop_479_480 top479 top480 {l}
Rbot_479_480 bot479 bot480 {r}
Lbot_479_480 bot479 bot480 {l}
Rtop_479_509 top479 top509 {r}
Ltop_479_509 top479 top509 {l}
Rbot_479_509 bot479 bot509 {r}
Lbot_479_509 bot479 bot509 {l}
C479 top479 bot479 {c}
Rtop_480_510 top480 top510 {r}
Ltop_480_510 top480 top510 {l}
Rbot_480_510 bot480 bot510 {r}
Lbot_480_510 bot480 bot510 {l}
C480 top480 bot480 {c}
Rtop_481_482 top481 top482 {r}
Ltop_481_482 top481 top482 {l}
Rbot_481_482 bot481 bot482 {r}
Lbot_481_482 bot481 bot482 {l}
Rtop_481_511 top481 top511 {r}
Ltop_481_511 top481 top511 {l}
Rbot_481_511 bot481 bot511 {r}
Lbot_481_511 bot481 bot511 {l}
C481 top481 bot481 {c}
Rtop_482_483 top482 top483 {r}
Ltop_482_483 top482 top483 {l}
Rbot_482_483 bot482 bot483 {r}
Lbot_482_483 bot482 bot483 {l}
Rtop_482_512 top482 top512 {r}
Ltop_482_512 top482 top512 {l}
Rbot_482_512 bot482 bot512 {r}
Lbot_482_512 bot482 bot512 {l}
C482 top482 bot482 {c}
Rtop_483_484 top483 top484 {r}
Ltop_483_484 top483 top484 {l}
Rbot_483_484 bot483 bot484 {r}
Lbot_483_484 bot483 bot484 {l}
Rtop_483_513 top483 top513 {r}
Ltop_483_513 top483 top513 {l}
Rbot_483_513 bot483 bot513 {r}
Lbot_483_513 bot483 bot513 {l}
C483 top483 bot483 {c}
Rtop_484_485 top484 top485 {r}
Ltop_484_485 top484 top485 {l}
Rbot_484_485 bot484 bot485 {r}
Lbot_484_485 bot484 bot485 {l}
Rtop_484_514 top484 top514 {r}
Ltop_484_514 top484 top514 {l}
Rbot_484_514 bot484 bot514 {r}
Lbot_484_514 bot484 bot514 {l}
C484 top484 bot484 {c}
Rtop_485_486 top485 top486 {r}
Ltop_485_486 top485 top486 {l}
Rbot_485_486 bot485 bot486 {r}
Lbot_485_486 bot485 bot486 {l}
Rtop_485_515 top485 top515 {r}
Ltop_485_515 top485 top515 {l}
Rbot_485_515 bot485 bot515 {r}
Lbot_485_515 bot485 bot515 {l}
C485 top485 bot485 {c}
Rtop_486_487 top486 top487 {r}
Ltop_486_487 top486 top487 {l}
Rbot_486_487 bot486 bot487 {r}
Lbot_486_487 bot486 bot487 {l}
Rtop_486_516 top486 top516 {r}
Ltop_486_516 top486 top516 {l}
Rbot_486_516 bot486 bot516 {r}
Lbot_486_516 bot486 bot516 {l}
C486 top486 bot486 {c}
Rtop_487_488 top487 top488 {r}
Ltop_487_488 top487 top488 {l}
Rbot_487_488 bot487 bot488 {r}
Lbot_487_488 bot487 bot488 {l}
Rtop_487_517 top487 top517 {r}
Ltop_487_517 top487 top517 {l}
Rbot_487_517 bot487 bot517 {r}
Lbot_487_517 bot487 bot517 {l}
C487 top487 bot487 {c}
Rtop_488_489 top488 top489 {r}
Ltop_488_489 top488 top489 {l}
Rbot_488_489 bot488 bot489 {r}
Lbot_488_489 bot488 bot489 {l}
Rtop_488_518 top488 top518 {r}
Ltop_488_518 top488 top518 {l}
Rbot_488_518 bot488 bot518 {r}
Lbot_488_518 bot488 bot518 {l}
C488 top488 bot488 {c}
Rtop_489_490 top489 top490 {r}
Ltop_489_490 top489 top490 {l}
Rbot_489_490 bot489 bot490 {r}
Lbot_489_490 bot489 bot490 {l}
Rtop_489_519 top489 top519 {r}
Ltop_489_519 top489 top519 {l}
Rbot_489_519 bot489 bot519 {r}
Lbot_489_519 bot489 bot519 {l}
C489 top489 bot489 {c}
Rtop_490_491 top490 top491 {r}
Ltop_490_491 top490 top491 {l}
Rbot_490_491 bot490 bot491 {r}
Lbot_490_491 bot490 bot491 {l}
Rtop_490_520 top490 top520 {r}
Ltop_490_520 top490 top520 {l}
Rbot_490_520 bot490 bot520 {r}
Lbot_490_520 bot490 bot520 {l}
C490 top490 bot490 {c}
Rtop_491_492 top491 top492 {r}
Ltop_491_492 top491 top492 {l}
Rbot_491_492 bot491 bot492 {r}
Lbot_491_492 bot491 bot492 {l}
Rtop_491_521 top491 top521 {r}
Ltop_491_521 top491 top521 {l}
Rbot_491_521 bot491 bot521 {r}
Lbot_491_521 bot491 bot521 {l}
C491 top491 bot491 {c}
Rtop_492_493 top492 top493 {r}
Ltop_492_493 top492 top493 {l}
Rbot_492_493 bot492 bot493 {r}
Lbot_492_493 bot492 bot493 {l}
Rtop_492_522 top492 top522 {r}
Ltop_492_522 top492 top522 {l}
Rbot_492_522 bot492 bot522 {r}
Lbot_492_522 bot492 bot522 {l}
C492 top492 bot492 {c}
Rtop_493_494 top493 top494 {r}
Ltop_493_494 top493 top494 {l}
Rbot_493_494 bot493 bot494 {r}
Lbot_493_494 bot493 bot494 {l}
Rtop_493_523 top493 top523 {r}
Ltop_493_523 top493 top523 {l}
Rbot_493_523 bot493 bot523 {r}
Lbot_493_523 bot493 bot523 {l}
C493 top493 bot493 {c}
Rtop_494_495 top494 top495 {r}
Ltop_494_495 top494 top495 {l}
Rbot_494_495 bot494 bot495 {r}
Lbot_494_495 bot494 bot495 {l}
Rtop_494_524 top494 top524 {r}
Ltop_494_524 top494 top524 {l}
Rbot_494_524 bot494 bot524 {r}
Lbot_494_524 bot494 bot524 {l}
C494 top494 bot494 {c}
Rtop_495_496 top495 top496 {r}
Ltop_495_496 top495 top496 {l}
Rbot_495_496 bot495 bot496 {r}
Lbot_495_496 bot495 bot496 {l}
Rtop_495_525 top495 top525 {r}
Ltop_495_525 top495 top525 {l}
Rbot_495_525 bot495 bot525 {r}
Lbot_495_525 bot495 bot525 {l}
C495 top495 bot495 {c}
Rtop_496_497 top496 top497 {r}
Ltop_496_497 top496 top497 {l}
Rbot_496_497 bot496 bot497 {r}
Lbot_496_497 bot496 bot497 {l}
Rtop_496_526 top496 top526 {r}
Ltop_496_526 top496 top526 {l}
Rbot_496_526 bot496 bot526 {r}
Lbot_496_526 bot496 bot526 {l}
C496 top496 bot496 {c}
Rtop_497_498 top497 top498 {r}
Ltop_497_498 top497 top498 {l}
Rbot_497_498 bot497 bot498 {r}
Lbot_497_498 bot497 bot498 {l}
Rtop_497_527 top497 top527 {r}
Ltop_497_527 top497 top527 {l}
Rbot_497_527 bot497 bot527 {r}
Lbot_497_527 bot497 bot527 {l}
C497 top497 bot497 {c}
Rtop_498_499 top498 top499 {r}
Ltop_498_499 top498 top499 {l}
Rbot_498_499 bot498 bot499 {r}
Lbot_498_499 bot498 bot499 {l}
Rtop_498_528 top498 top528 {r}
Ltop_498_528 top498 top528 {l}
Rbot_498_528 bot498 bot528 {r}
Lbot_498_528 bot498 bot528 {l}
C498 top498 bot498 {c}
Rtop_499_500 top499 top500 {r}
Ltop_499_500 top499 top500 {l}
Rbot_499_500 bot499 bot500 {r}
Lbot_499_500 bot499 bot500 {l}
Rtop_499_529 top499 top529 {r}
Ltop_499_529 top499 top529 {l}
Rbot_499_529 bot499 bot529 {r}
Lbot_499_529 bot499 bot529 {l}
C499 top499 bot499 {c}
Rtop_500_501 top500 top501 {r}
Ltop_500_501 top500 top501 {l}
Rbot_500_501 bot500 bot501 {r}
Lbot_500_501 bot500 bot501 {l}
Rtop_500_530 top500 top530 {r}
Ltop_500_530 top500 top530 {l}
Rbot_500_530 bot500 bot530 {r}
Lbot_500_530 bot500 bot530 {l}
C500 top500 bot500 {c}
Rtop_501_502 top501 top502 {r}
Ltop_501_502 top501 top502 {l}
Rbot_501_502 bot501 bot502 {r}
Lbot_501_502 bot501 bot502 {l}
Rtop_501_531 top501 top531 {r}
Ltop_501_531 top501 top531 {l}
Rbot_501_531 bot501 bot531 {r}
Lbot_501_531 bot501 bot531 {l}
C501 top501 bot501 {c}
Rtop_502_503 top502 top503 {r}
Ltop_502_503 top502 top503 {l}
Rbot_502_503 bot502 bot503 {r}
Lbot_502_503 bot502 bot503 {l}
Rtop_502_532 top502 top532 {r}
Ltop_502_532 top502 top532 {l}
Rbot_502_532 bot502 bot532 {r}
Lbot_502_532 bot502 bot532 {l}
C502 top502 bot502 {c}
Rtop_503_504 top503 top504 {r}
Ltop_503_504 top503 top504 {l}
Rbot_503_504 bot503 bot504 {r}
Lbot_503_504 bot503 bot504 {l}
Rtop_503_533 top503 top533 {r}
Ltop_503_533 top503 top533 {l}
Rbot_503_533 bot503 bot533 {r}
Lbot_503_533 bot503 bot533 {l}
C503 top503 bot503 {c}
Rtop_504_505 top504 top505 {r}
Ltop_504_505 top504 top505 {l}
Rbot_504_505 bot504 bot505 {r}
Lbot_504_505 bot504 bot505 {l}
Rtop_504_534 top504 top534 {r}
Ltop_504_534 top504 top534 {l}
Rbot_504_534 bot504 bot534 {r}
Lbot_504_534 bot504 bot534 {l}
C504 top504 bot504 {c}
Rtop_505_506 top505 top506 {r}
Ltop_505_506 top505 top506 {l}
Rbot_505_506 bot505 bot506 {r}
Lbot_505_506 bot505 bot506 {l}
Rtop_505_535 top505 top535 {r}
Ltop_505_535 top505 top535 {l}
Rbot_505_535 bot505 bot535 {r}
Lbot_505_535 bot505 bot535 {l}
C505 top505 bot505 {c}
Rtop_506_507 top506 top507 {r}
Ltop_506_507 top506 top507 {l}
Rbot_506_507 bot506 bot507 {r}
Lbot_506_507 bot506 bot507 {l}
Rtop_506_536 top506 top536 {r}
Ltop_506_536 top506 top536 {l}
Rbot_506_536 bot506 bot536 {r}
Lbot_506_536 bot506 bot536 {l}
C506 top506 bot506 {c}
Rtop_507_508 top507 top508 {r}
Ltop_507_508 top507 top508 {l}
Rbot_507_508 bot507 bot508 {r}
Lbot_507_508 bot507 bot508 {l}
Rtop_507_537 top507 top537 {r}
Ltop_507_537 top507 top537 {l}
Rbot_507_537 bot507 bot537 {r}
Lbot_507_537 bot507 bot537 {l}
C507 top507 bot507 {c}
Rtop_508_509 top508 top509 {r}
Ltop_508_509 top508 top509 {l}
Rbot_508_509 bot508 bot509 {r}
Lbot_508_509 bot508 bot509 {l}
Rtop_508_538 top508 top538 {r}
Ltop_508_538 top508 top538 {l}
Rbot_508_538 bot508 bot538 {r}
Lbot_508_538 bot508 bot538 {l}
C508 top508 bot508 {c}
Rtop_509_510 top509 top510 {r}
Ltop_509_510 top509 top510 {l}
Rbot_509_510 bot509 bot510 {r}
Lbot_509_510 bot509 bot510 {l}
Rtop_509_539 top509 top539 {r}
Ltop_509_539 top509 top539 {l}
Rbot_509_539 bot509 bot539 {r}
Lbot_509_539 bot509 bot539 {l}
C509 top509 bot509 {c}
Rtop_510_540 top510 top540 {r}
Ltop_510_540 top510 top540 {l}
Rbot_510_540 bot510 bot540 {r}
Lbot_510_540 bot510 bot540 {l}
C510 top510 bot510 {c}
Rtop_511_512 top511 top512 {r}
Ltop_511_512 top511 top512 {l}
Rbot_511_512 bot511 bot512 {r}
Lbot_511_512 bot511 bot512 {l}
Rtop_511_541 top511 top541 {r}
Ltop_511_541 top511 top541 {l}
Rbot_511_541 bot511 bot541 {r}
Lbot_511_541 bot511 bot541 {l}
C511 top511 bot511 {c}
Rtop_512_513 top512 top513 {r}
Ltop_512_513 top512 top513 {l}
Rbot_512_513 bot512 bot513 {r}
Lbot_512_513 bot512 bot513 {l}
Rtop_512_542 top512 top542 {r}
Ltop_512_542 top512 top542 {l}
Rbot_512_542 bot512 bot542 {r}
Lbot_512_542 bot512 bot542 {l}
C512 top512 bot512 {c}
Rtop_513_514 top513 top514 {r}
Ltop_513_514 top513 top514 {l}
Rbot_513_514 bot513 bot514 {r}
Lbot_513_514 bot513 bot514 {l}
Rtop_513_543 top513 top543 {r}
Ltop_513_543 top513 top543 {l}
Rbot_513_543 bot513 bot543 {r}
Lbot_513_543 bot513 bot543 {l}
C513 top513 bot513 {c}
Rtop_514_515 top514 top515 {r}
Ltop_514_515 top514 top515 {l}
Rbot_514_515 bot514 bot515 {r}
Lbot_514_515 bot514 bot515 {l}
Rtop_514_544 top514 top544 {r}
Ltop_514_544 top514 top544 {l}
Rbot_514_544 bot514 bot544 {r}
Lbot_514_544 bot514 bot544 {l}
C514 top514 bot514 {c}
Rtop_515_516 top515 top516 {r}
Ltop_515_516 top515 top516 {l}
Rbot_515_516 bot515 bot516 {r}
Lbot_515_516 bot515 bot516 {l}
Rtop_515_545 top515 top545 {r}
Ltop_515_545 top515 top545 {l}
Rbot_515_545 bot515 bot545 {r}
Lbot_515_545 bot515 bot545 {l}
C515 top515 bot515 {c}
Rtop_516_517 top516 top517 {r}
Ltop_516_517 top516 top517 {l}
Rbot_516_517 bot516 bot517 {r}
Lbot_516_517 bot516 bot517 {l}
Rtop_516_546 top516 top546 {r}
Ltop_516_546 top516 top546 {l}
Rbot_516_546 bot516 bot546 {r}
Lbot_516_546 bot516 bot546 {l}
C516 top516 bot516 {c}
Rtop_517_518 top517 top518 {r}
Ltop_517_518 top517 top518 {l}
Rbot_517_518 bot517 bot518 {r}
Lbot_517_518 bot517 bot518 {l}
Rtop_517_547 top517 top547 {r}
Ltop_517_547 top517 top547 {l}
Rbot_517_547 bot517 bot547 {r}
Lbot_517_547 bot517 bot547 {l}
C517 top517 bot517 {c}
Rtop_518_519 top518 top519 {r}
Ltop_518_519 top518 top519 {l}
Rbot_518_519 bot518 bot519 {r}
Lbot_518_519 bot518 bot519 {l}
Rtop_518_548 top518 top548 {r}
Ltop_518_548 top518 top548 {l}
Rbot_518_548 bot518 bot548 {r}
Lbot_518_548 bot518 bot548 {l}
C518 top518 bot518 {c}
Rtop_519_520 top519 top520 {r}
Ltop_519_520 top519 top520 {l}
Rbot_519_520 bot519 bot520 {r}
Lbot_519_520 bot519 bot520 {l}
Rtop_519_549 top519 top549 {r}
Ltop_519_549 top519 top549 {l}
Rbot_519_549 bot519 bot549 {r}
Lbot_519_549 bot519 bot549 {l}
C519 top519 bot519 {c}
Rtop_520_521 top520 top521 {r}
Ltop_520_521 top520 top521 {l}
Rbot_520_521 bot520 bot521 {r}
Lbot_520_521 bot520 bot521 {l}
Rtop_520_550 top520 top550 {r}
Ltop_520_550 top520 top550 {l}
Rbot_520_550 bot520 bot550 {r}
Lbot_520_550 bot520 bot550 {l}
C520 top520 bot520 {c}
Rtop_521_522 top521 top522 {r}
Ltop_521_522 top521 top522 {l}
Rbot_521_522 bot521 bot522 {r}
Lbot_521_522 bot521 bot522 {l}
Rtop_521_551 top521 top551 {r}
Ltop_521_551 top521 top551 {l}
Rbot_521_551 bot521 bot551 {r}
Lbot_521_551 bot521 bot551 {l}
C521 top521 bot521 {c}
Rtop_522_523 top522 top523 {r}
Ltop_522_523 top522 top523 {l}
Rbot_522_523 bot522 bot523 {r}
Lbot_522_523 bot522 bot523 {l}
Rtop_522_552 top522 top552 {r}
Ltop_522_552 top522 top552 {l}
Rbot_522_552 bot522 bot552 {r}
Lbot_522_552 bot522 bot552 {l}
C522 top522 bot522 {c}
Rtop_523_524 top523 top524 {r}
Ltop_523_524 top523 top524 {l}
Rbot_523_524 bot523 bot524 {r}
Lbot_523_524 bot523 bot524 {l}
Rtop_523_553 top523 top553 {r}
Ltop_523_553 top523 top553 {l}
Rbot_523_553 bot523 bot553 {r}
Lbot_523_553 bot523 bot553 {l}
C523 top523 bot523 {c}
Rtop_524_525 top524 top525 {r}
Ltop_524_525 top524 top525 {l}
Rbot_524_525 bot524 bot525 {r}
Lbot_524_525 bot524 bot525 {l}
Rtop_524_554 top524 top554 {r}
Ltop_524_554 top524 top554 {l}
Rbot_524_554 bot524 bot554 {r}
Lbot_524_554 bot524 bot554 {l}
C524 top524 bot524 {c}
Rtop_525_526 top525 top526 {r}
Ltop_525_526 top525 top526 {l}
Rbot_525_526 bot525 bot526 {r}
Lbot_525_526 bot525 bot526 {l}
Rtop_525_555 top525 top555 {r}
Ltop_525_555 top525 top555 {l}
Rbot_525_555 bot525 bot555 {r}
Lbot_525_555 bot525 bot555 {l}
C525 top525 bot525 {c}
Rtop_526_527 top526 top527 {r}
Ltop_526_527 top526 top527 {l}
Rbot_526_527 bot526 bot527 {r}
Lbot_526_527 bot526 bot527 {l}
Rtop_526_556 top526 top556 {r}
Ltop_526_556 top526 top556 {l}
Rbot_526_556 bot526 bot556 {r}
Lbot_526_556 bot526 bot556 {l}
C526 top526 bot526 {c}
Rtop_527_528 top527 top528 {r}
Ltop_527_528 top527 top528 {l}
Rbot_527_528 bot527 bot528 {r}
Lbot_527_528 bot527 bot528 {l}
Rtop_527_557 top527 top557 {r}
Ltop_527_557 top527 top557 {l}
Rbot_527_557 bot527 bot557 {r}
Lbot_527_557 bot527 bot557 {l}
C527 top527 bot527 {c}
Rtop_528_529 top528 top529 {r}
Ltop_528_529 top528 top529 {l}
Rbot_528_529 bot528 bot529 {r}
Lbot_528_529 bot528 bot529 {l}
Rtop_528_558 top528 top558 {r}
Ltop_528_558 top528 top558 {l}
Rbot_528_558 bot528 bot558 {r}
Lbot_528_558 bot528 bot558 {l}
C528 top528 bot528 {c}
Rtop_529_530 top529 top530 {r}
Ltop_529_530 top529 top530 {l}
Rbot_529_530 bot529 bot530 {r}
Lbot_529_530 bot529 bot530 {l}
Rtop_529_559 top529 top559 {r}
Ltop_529_559 top529 top559 {l}
Rbot_529_559 bot529 bot559 {r}
Lbot_529_559 bot529 bot559 {l}
C529 top529 bot529 {c}
Rtop_530_531 top530 top531 {r}
Ltop_530_531 top530 top531 {l}
Rbot_530_531 bot530 bot531 {r}
Lbot_530_531 bot530 bot531 {l}
Rtop_530_560 top530 top560 {r}
Ltop_530_560 top530 top560 {l}
Rbot_530_560 bot530 bot560 {r}
Lbot_530_560 bot530 bot560 {l}
C530 top530 bot530 {c}
Rtop_531_532 top531 top532 {r}
Ltop_531_532 top531 top532 {l}
Rbot_531_532 bot531 bot532 {r}
Lbot_531_532 bot531 bot532 {l}
Rtop_531_561 top531 top561 {r}
Ltop_531_561 top531 top561 {l}
Rbot_531_561 bot531 bot561 {r}
Lbot_531_561 bot531 bot561 {l}
C531 top531 bot531 {c}
Rtop_532_533 top532 top533 {r}
Ltop_532_533 top532 top533 {l}
Rbot_532_533 bot532 bot533 {r}
Lbot_532_533 bot532 bot533 {l}
Rtop_532_562 top532 top562 {r}
Ltop_532_562 top532 top562 {l}
Rbot_532_562 bot532 bot562 {r}
Lbot_532_562 bot532 bot562 {l}
C532 top532 bot532 {c}
Rtop_533_534 top533 top534 {r}
Ltop_533_534 top533 top534 {l}
Rbot_533_534 bot533 bot534 {r}
Lbot_533_534 bot533 bot534 {l}
Rtop_533_563 top533 top563 {r}
Ltop_533_563 top533 top563 {l}
Rbot_533_563 bot533 bot563 {r}
Lbot_533_563 bot533 bot563 {l}
C533 top533 bot533 {c}
Rtop_534_535 top534 top535 {r}
Ltop_534_535 top534 top535 {l}
Rbot_534_535 bot534 bot535 {r}
Lbot_534_535 bot534 bot535 {l}
Rtop_534_564 top534 top564 {r}
Ltop_534_564 top534 top564 {l}
Rbot_534_564 bot534 bot564 {r}
Lbot_534_564 bot534 bot564 {l}
C534 top534 bot534 {c}
Rtop_535_536 top535 top536 {r}
Ltop_535_536 top535 top536 {l}
Rbot_535_536 bot535 bot536 {r}
Lbot_535_536 bot535 bot536 {l}
Rtop_535_565 top535 top565 {r}
Ltop_535_565 top535 top565 {l}
Rbot_535_565 bot535 bot565 {r}
Lbot_535_565 bot535 bot565 {l}
C535 top535 bot535 {c}
Rtop_536_537 top536 top537 {r}
Ltop_536_537 top536 top537 {l}
Rbot_536_537 bot536 bot537 {r}
Lbot_536_537 bot536 bot537 {l}
Rtop_536_566 top536 top566 {r}
Ltop_536_566 top536 top566 {l}
Rbot_536_566 bot536 bot566 {r}
Lbot_536_566 bot536 bot566 {l}
C536 top536 bot536 {c}
Rtop_537_538 top537 top538 {r}
Ltop_537_538 top537 top538 {l}
Rbot_537_538 bot537 bot538 {r}
Lbot_537_538 bot537 bot538 {l}
Rtop_537_567 top537 top567 {r}
Ltop_537_567 top537 top567 {l}
Rbot_537_567 bot537 bot567 {r}
Lbot_537_567 bot537 bot567 {l}
C537 top537 bot537 {c}
Rtop_538_539 top538 top539 {r}
Ltop_538_539 top538 top539 {l}
Rbot_538_539 bot538 bot539 {r}
Lbot_538_539 bot538 bot539 {l}
Rtop_538_568 top538 top568 {r}
Ltop_538_568 top538 top568 {l}
Rbot_538_568 bot538 bot568 {r}
Lbot_538_568 bot538 bot568 {l}
C538 top538 bot538 {c}
Rtop_539_540 top539 top540 {r}
Ltop_539_540 top539 top540 {l}
Rbot_539_540 bot539 bot540 {r}
Lbot_539_540 bot539 bot540 {l}
Rtop_539_569 top539 top569 {r}
Ltop_539_569 top539 top569 {l}
Rbot_539_569 bot539 bot569 {r}
Lbot_539_569 bot539 bot569 {l}
C539 top539 bot539 {c}
Rtop_540_570 top540 top570 {r}
Ltop_540_570 top540 top570 {l}
Rbot_540_570 bot540 bot570 {r}
Lbot_540_570 bot540 bot570 {l}
C540 top540 bot540 {c}
Rtop_541_542 top541 top542 {r}
Ltop_541_542 top541 top542 {l}
Rbot_541_542 bot541 bot542 {r}
Lbot_541_542 bot541 bot542 {l}
Rtop_541_571 top541 top571 {r}
Ltop_541_571 top541 top571 {l}
Rbot_541_571 bot541 bot571 {r}
Lbot_541_571 bot541 bot571 {l}
C541 top541 bot541 {c}
Rtop_542_543 top542 top543 {r}
Ltop_542_543 top542 top543 {l}
Rbot_542_543 bot542 bot543 {r}
Lbot_542_543 bot542 bot543 {l}
Rtop_542_572 top542 top572 {r}
Ltop_542_572 top542 top572 {l}
Rbot_542_572 bot542 bot572 {r}
Lbot_542_572 bot542 bot572 {l}
C542 top542 bot542 {c}
Rtop_543_544 top543 top544 {r}
Ltop_543_544 top543 top544 {l}
Rbot_543_544 bot543 bot544 {r}
Lbot_543_544 bot543 bot544 {l}
Rtop_543_573 top543 top573 {r}
Ltop_543_573 top543 top573 {l}
Rbot_543_573 bot543 bot573 {r}
Lbot_543_573 bot543 bot573 {l}
C543 top543 bot543 {c}
Rtop_544_545 top544 top545 {r}
Ltop_544_545 top544 top545 {l}
Rbot_544_545 bot544 bot545 {r}
Lbot_544_545 bot544 bot545 {l}
Rtop_544_574 top544 top574 {r}
Ltop_544_574 top544 top574 {l}
Rbot_544_574 bot544 bot574 {r}
Lbot_544_574 bot544 bot574 {l}
C544 top544 bot544 {c}
Rtop_545_546 top545 top546 {r}
Ltop_545_546 top545 top546 {l}
Rbot_545_546 bot545 bot546 {r}
Lbot_545_546 bot545 bot546 {l}
Rtop_545_575 top545 top575 {r}
Ltop_545_575 top545 top575 {l}
Rbot_545_575 bot545 bot575 {r}
Lbot_545_575 bot545 bot575 {l}
C545 top545 bot545 {c}
Rtop_546_547 top546 top547 {r}
Ltop_546_547 top546 top547 {l}
Rbot_546_547 bot546 bot547 {r}
Lbot_546_547 bot546 bot547 {l}
Rtop_546_576 top546 top576 {r}
Ltop_546_576 top546 top576 {l}
Rbot_546_576 bot546 bot576 {r}
Lbot_546_576 bot546 bot576 {l}
C546 top546 bot546 {c}
Rtop_547_548 top547 top548 {r}
Ltop_547_548 top547 top548 {l}
Rbot_547_548 bot547 bot548 {r}
Lbot_547_548 bot547 bot548 {l}
Rtop_547_577 top547 top577 {r}
Ltop_547_577 top547 top577 {l}
Rbot_547_577 bot547 bot577 {r}
Lbot_547_577 bot547 bot577 {l}
C547 top547 bot547 {c}
Rtop_548_549 top548 top549 {r}
Ltop_548_549 top548 top549 {l}
Rbot_548_549 bot548 bot549 {r}
Lbot_548_549 bot548 bot549 {l}
Rtop_548_578 top548 top578 {r}
Ltop_548_578 top548 top578 {l}
Rbot_548_578 bot548 bot578 {r}
Lbot_548_578 bot548 bot578 {l}
C548 top548 bot548 {c}
Rtop_549_550 top549 top550 {r}
Ltop_549_550 top549 top550 {l}
Rbot_549_550 bot549 bot550 {r}
Lbot_549_550 bot549 bot550 {l}
Rtop_549_579 top549 top579 {r}
Ltop_549_579 top549 top579 {l}
Rbot_549_579 bot549 bot579 {r}
Lbot_549_579 bot549 bot579 {l}
C549 top549 bot549 {c}
Rtop_550_551 top550 top551 {r}
Ltop_550_551 top550 top551 {l}
Rbot_550_551 bot550 bot551 {r}
Lbot_550_551 bot550 bot551 {l}
Rtop_550_580 top550 top580 {r}
Ltop_550_580 top550 top580 {l}
Rbot_550_580 bot550 bot580 {r}
Lbot_550_580 bot550 bot580 {l}
C550 top550 bot550 {c}
Rtop_551_552 top551 top552 {r}
Ltop_551_552 top551 top552 {l}
Rbot_551_552 bot551 bot552 {r}
Lbot_551_552 bot551 bot552 {l}
Rtop_551_581 top551 top581 {r}
Ltop_551_581 top551 top581 {l}
Rbot_551_581 bot551 bot581 {r}
Lbot_551_581 bot551 bot581 {l}
C551 top551 bot551 {c}
Rtop_552_553 top552 top553 {r}
Ltop_552_553 top552 top553 {l}
Rbot_552_553 bot552 bot553 {r}
Lbot_552_553 bot552 bot553 {l}
Rtop_552_582 top552 top582 {r}
Ltop_552_582 top552 top582 {l}
Rbot_552_582 bot552 bot582 {r}
Lbot_552_582 bot552 bot582 {l}
C552 top552 bot552 {c}
Rtop_553_554 top553 top554 {r}
Ltop_553_554 top553 top554 {l}
Rbot_553_554 bot553 bot554 {r}
Lbot_553_554 bot553 bot554 {l}
Rtop_553_583 top553 top583 {r}
Ltop_553_583 top553 top583 {l}
Rbot_553_583 bot553 bot583 {r}
Lbot_553_583 bot553 bot583 {l}
C553 top553 bot553 {c}
Rtop_554_555 top554 top555 {r}
Ltop_554_555 top554 top555 {l}
Rbot_554_555 bot554 bot555 {r}
Lbot_554_555 bot554 bot555 {l}
Rtop_554_584 top554 top584 {r}
Ltop_554_584 top554 top584 {l}
Rbot_554_584 bot554 bot584 {r}
Lbot_554_584 bot554 bot584 {l}
C554 top554 bot554 {c}
Rtop_555_556 top555 top556 {r}
Ltop_555_556 top555 top556 {l}
Rbot_555_556 bot555 bot556 {r}
Lbot_555_556 bot555 bot556 {l}
Rtop_555_585 top555 top585 {r}
Ltop_555_585 top555 top585 {l}
Rbot_555_585 bot555 bot585 {r}
Lbot_555_585 bot555 bot585 {l}
C555 top555 bot555 {c}
Rtop_556_557 top556 top557 {r}
Ltop_556_557 top556 top557 {l}
Rbot_556_557 bot556 bot557 {r}
Lbot_556_557 bot556 bot557 {l}
Rtop_556_586 top556 top586 {r}
Ltop_556_586 top556 top586 {l}
Rbot_556_586 bot556 bot586 {r}
Lbot_556_586 bot556 bot586 {l}
C556 top556 bot556 {c}
Rtop_557_558 top557 top558 {r}
Ltop_557_558 top557 top558 {l}
Rbot_557_558 bot557 bot558 {r}
Lbot_557_558 bot557 bot558 {l}
Rtop_557_587 top557 top587 {r}
Ltop_557_587 top557 top587 {l}
Rbot_557_587 bot557 bot587 {r}
Lbot_557_587 bot557 bot587 {l}
C557 top557 bot557 {c}
Rtop_558_559 top558 top559 {r}
Ltop_558_559 top558 top559 {l}
Rbot_558_559 bot558 bot559 {r}
Lbot_558_559 bot558 bot559 {l}
Rtop_558_588 top558 top588 {r}
Ltop_558_588 top558 top588 {l}
Rbot_558_588 bot558 bot588 {r}
Lbot_558_588 bot558 bot588 {l}
C558 top558 bot558 {c}
Rtop_559_560 top559 top560 {r}
Ltop_559_560 top559 top560 {l}
Rbot_559_560 bot559 bot560 {r}
Lbot_559_560 bot559 bot560 {l}
Rtop_559_589 top559 top589 {r}
Ltop_559_589 top559 top589 {l}
Rbot_559_589 bot559 bot589 {r}
Lbot_559_589 bot559 bot589 {l}
C559 top559 bot559 {c}
Rtop_560_561 top560 top561 {r}
Ltop_560_561 top560 top561 {l}
Rbot_560_561 bot560 bot561 {r}
Lbot_560_561 bot560 bot561 {l}
Rtop_560_590 top560 top590 {r}
Ltop_560_590 top560 top590 {l}
Rbot_560_590 bot560 bot590 {r}
Lbot_560_590 bot560 bot590 {l}
C560 top560 bot560 {c}
Rtop_561_562 top561 top562 {r}
Ltop_561_562 top561 top562 {l}
Rbot_561_562 bot561 bot562 {r}
Lbot_561_562 bot561 bot562 {l}
Rtop_561_591 top561 top591 {r}
Ltop_561_591 top561 top591 {l}
Rbot_561_591 bot561 bot591 {r}
Lbot_561_591 bot561 bot591 {l}
C561 top561 bot561 {c}
Rtop_562_563 top562 top563 {r}
Ltop_562_563 top562 top563 {l}
Rbot_562_563 bot562 bot563 {r}
Lbot_562_563 bot562 bot563 {l}
Rtop_562_592 top562 top592 {r}
Ltop_562_592 top562 top592 {l}
Rbot_562_592 bot562 bot592 {r}
Lbot_562_592 bot562 bot592 {l}
C562 top562 bot562 {c}
Rtop_563_564 top563 top564 {r}
Ltop_563_564 top563 top564 {l}
Rbot_563_564 bot563 bot564 {r}
Lbot_563_564 bot563 bot564 {l}
Rtop_563_593 top563 top593 {r}
Ltop_563_593 top563 top593 {l}
Rbot_563_593 bot563 bot593 {r}
Lbot_563_593 bot563 bot593 {l}
C563 top563 bot563 {c}
Rtop_564_565 top564 top565 {r}
Ltop_564_565 top564 top565 {l}
Rbot_564_565 bot564 bot565 {r}
Lbot_564_565 bot564 bot565 {l}
Rtop_564_594 top564 top594 {r}
Ltop_564_594 top564 top594 {l}
Rbot_564_594 bot564 bot594 {r}
Lbot_564_594 bot564 bot594 {l}
C564 top564 bot564 {c}
Rtop_565_566 top565 top566 {r}
Ltop_565_566 top565 top566 {l}
Rbot_565_566 bot565 bot566 {r}
Lbot_565_566 bot565 bot566 {l}
Rtop_565_595 top565 top595 {r}
Ltop_565_595 top565 top595 {l}
Rbot_565_595 bot565 bot595 {r}
Lbot_565_595 bot565 bot595 {l}
C565 top565 bot565 {c}
Rtop_566_567 top566 top567 {r}
Ltop_566_567 top566 top567 {l}
Rbot_566_567 bot566 bot567 {r}
Lbot_566_567 bot566 bot567 {l}
Rtop_566_596 top566 top596 {r}
Ltop_566_596 top566 top596 {l}
Rbot_566_596 bot566 bot596 {r}
Lbot_566_596 bot566 bot596 {l}
C566 top566 bot566 {c}
Rtop_567_568 top567 top568 {r}
Ltop_567_568 top567 top568 {l}
Rbot_567_568 bot567 bot568 {r}
Lbot_567_568 bot567 bot568 {l}
Rtop_567_597 top567 top597 {r}
Ltop_567_597 top567 top597 {l}
Rbot_567_597 bot567 bot597 {r}
Lbot_567_597 bot567 bot597 {l}
C567 top567 bot567 {c}
Rtop_568_569 top568 top569 {r}
Ltop_568_569 top568 top569 {l}
Rbot_568_569 bot568 bot569 {r}
Lbot_568_569 bot568 bot569 {l}
Rtop_568_598 top568 top598 {r}
Ltop_568_598 top568 top598 {l}
Rbot_568_598 bot568 bot598 {r}
Lbot_568_598 bot568 bot598 {l}
C568 top568 bot568 {c}
Rtop_569_570 top569 top570 {r}
Ltop_569_570 top569 top570 {l}
Rbot_569_570 bot569 bot570 {r}
Lbot_569_570 bot569 bot570 {l}
Rtop_569_599 top569 top599 {r}
Ltop_569_599 top569 top599 {l}
Rbot_569_599 bot569 bot599 {r}
Lbot_569_599 bot569 bot599 {l}
C569 top569 bot569 {c}
Rtop_570_600 top570 top600 {r}
Ltop_570_600 top570 top600 {l}
Rbot_570_600 bot570 bot600 {r}
Lbot_570_600 bot570 bot600 {l}
C570 top570 bot570 {c}
Rtop_571_572 top571 top572 {r}
Ltop_571_572 top571 top572 {l}
Rbot_571_572 bot571 bot572 {r}
Lbot_571_572 bot571 bot572 {l}
Rtop_571_601 top571 top601 {r}
Ltop_571_601 top571 top601 {l}
Rbot_571_601 bot571 bot601 {r}
Lbot_571_601 bot571 bot601 {l}
C571 top571 bot571 {c}
Rtop_572_573 top572 top573 {r}
Ltop_572_573 top572 top573 {l}
Rbot_572_573 bot572 bot573 {r}
Lbot_572_573 bot572 bot573 {l}
Rtop_572_602 top572 top602 {r}
Ltop_572_602 top572 top602 {l}
Rbot_572_602 bot572 bot602 {r}
Lbot_572_602 bot572 bot602 {l}
C572 top572 bot572 {c}
Rtop_573_574 top573 top574 {r}
Ltop_573_574 top573 top574 {l}
Rbot_573_574 bot573 bot574 {r}
Lbot_573_574 bot573 bot574 {l}
Rtop_573_603 top573 top603 {r}
Ltop_573_603 top573 top603 {l}
Rbot_573_603 bot573 bot603 {r}
Lbot_573_603 bot573 bot603 {l}
C573 top573 bot573 {c}
Rtop_574_575 top574 top575 {r}
Ltop_574_575 top574 top575 {l}
Rbot_574_575 bot574 bot575 {r}
Lbot_574_575 bot574 bot575 {l}
Rtop_574_604 top574 top604 {r}
Ltop_574_604 top574 top604 {l}
Rbot_574_604 bot574 bot604 {r}
Lbot_574_604 bot574 bot604 {l}
C574 top574 bot574 {c}
Rtop_575_576 top575 top576 {r}
Ltop_575_576 top575 top576 {l}
Rbot_575_576 bot575 bot576 {r}
Lbot_575_576 bot575 bot576 {l}
Rtop_575_605 top575 top605 {r}
Ltop_575_605 top575 top605 {l}
Rbot_575_605 bot575 bot605 {r}
Lbot_575_605 bot575 bot605 {l}
C575 top575 bot575 {c}
Rtop_576_577 top576 top577 {r}
Ltop_576_577 top576 top577 {l}
Rbot_576_577 bot576 bot577 {r}
Lbot_576_577 bot576 bot577 {l}
Rtop_576_606 top576 top606 {r}
Ltop_576_606 top576 top606 {l}
Rbot_576_606 bot576 bot606 {r}
Lbot_576_606 bot576 bot606 {l}
C576 top576 bot576 {c}
Rtop_577_578 top577 top578 {r}
Ltop_577_578 top577 top578 {l}
Rbot_577_578 bot577 bot578 {r}
Lbot_577_578 bot577 bot578 {l}
Rtop_577_607 top577 top607 {r}
Ltop_577_607 top577 top607 {l}
Rbot_577_607 bot577 bot607 {r}
Lbot_577_607 bot577 bot607 {l}
C577 top577 bot577 {c}
Rtop_578_579 top578 top579 {r}
Ltop_578_579 top578 top579 {l}
Rbot_578_579 bot578 bot579 {r}
Lbot_578_579 bot578 bot579 {l}
Rtop_578_608 top578 top608 {r}
Ltop_578_608 top578 top608 {l}
Rbot_578_608 bot578 bot608 {r}
Lbot_578_608 bot578 bot608 {l}
C578 top578 bot578 {c}
Rtop_579_580 top579 top580 {r}
Ltop_579_580 top579 top580 {l}
Rbot_579_580 bot579 bot580 {r}
Lbot_579_580 bot579 bot580 {l}
Rtop_579_609 top579 top609 {r}
Ltop_579_609 top579 top609 {l}
Rbot_579_609 bot579 bot609 {r}
Lbot_579_609 bot579 bot609 {l}
C579 top579 bot579 {c}
Rtop_580_581 top580 top581 {r}
Ltop_580_581 top580 top581 {l}
Rbot_580_581 bot580 bot581 {r}
Lbot_580_581 bot580 bot581 {l}
Rtop_580_610 top580 top610 {r}
Ltop_580_610 top580 top610 {l}
Rbot_580_610 bot580 bot610 {r}
Lbot_580_610 bot580 bot610 {l}
C580 top580 bot580 {c}
Rtop_581_582 top581 top582 {r}
Ltop_581_582 top581 top582 {l}
Rbot_581_582 bot581 bot582 {r}
Lbot_581_582 bot581 bot582 {l}
Rtop_581_611 top581 top611 {r}
Ltop_581_611 top581 top611 {l}
Rbot_581_611 bot581 bot611 {r}
Lbot_581_611 bot581 bot611 {l}
C581 top581 bot581 {c}
Rtop_582_583 top582 top583 {r}
Ltop_582_583 top582 top583 {l}
Rbot_582_583 bot582 bot583 {r}
Lbot_582_583 bot582 bot583 {l}
Rtop_582_612 top582 top612 {r}
Ltop_582_612 top582 top612 {l}
Rbot_582_612 bot582 bot612 {r}
Lbot_582_612 bot582 bot612 {l}
C582 top582 bot582 {c}
Rtop_583_584 top583 top584 {r}
Ltop_583_584 top583 top584 {l}
Rbot_583_584 bot583 bot584 {r}
Lbot_583_584 bot583 bot584 {l}
Rtop_583_613 top583 top613 {r}
Ltop_583_613 top583 top613 {l}
Rbot_583_613 bot583 bot613 {r}
Lbot_583_613 bot583 bot613 {l}
C583 top583 bot583 {c}
Rtop_584_585 top584 top585 {r}
Ltop_584_585 top584 top585 {l}
Rbot_584_585 bot584 bot585 {r}
Lbot_584_585 bot584 bot585 {l}
Rtop_584_614 top584 top614 {r}
Ltop_584_614 top584 top614 {l}
Rbot_584_614 bot584 bot614 {r}
Lbot_584_614 bot584 bot614 {l}
C584 top584 bot584 {c}
Rtop_585_586 top585 top586 {r}
Ltop_585_586 top585 top586 {l}
Rbot_585_586 bot585 bot586 {r}
Lbot_585_586 bot585 bot586 {l}
Rtop_585_615 top585 top615 {r}
Ltop_585_615 top585 top615 {l}
Rbot_585_615 bot585 bot615 {r}
Lbot_585_615 bot585 bot615 {l}
C585 top585 bot585 {c}
Rtop_586_587 top586 top587 {r}
Ltop_586_587 top586 top587 {l}
Rbot_586_587 bot586 bot587 {r}
Lbot_586_587 bot586 bot587 {l}
Rtop_586_616 top586 top616 {r}
Ltop_586_616 top586 top616 {l}
Rbot_586_616 bot586 bot616 {r}
Lbot_586_616 bot586 bot616 {l}
C586 top586 bot586 {c}
Rtop_587_588 top587 top588 {r}
Ltop_587_588 top587 top588 {l}
Rbot_587_588 bot587 bot588 {r}
Lbot_587_588 bot587 bot588 {l}
Rtop_587_617 top587 top617 {r}
Ltop_587_617 top587 top617 {l}
Rbot_587_617 bot587 bot617 {r}
Lbot_587_617 bot587 bot617 {l}
C587 top587 bot587 {c}
Rtop_588_589 top588 top589 {r}
Ltop_588_589 top588 top589 {l}
Rbot_588_589 bot588 bot589 {r}
Lbot_588_589 bot588 bot589 {l}
Rtop_588_618 top588 top618 {r}
Ltop_588_618 top588 top618 {l}
Rbot_588_618 bot588 bot618 {r}
Lbot_588_618 bot588 bot618 {l}
C588 top588 bot588 {c}
Rtop_589_590 top589 top590 {r}
Ltop_589_590 top589 top590 {l}
Rbot_589_590 bot589 bot590 {r}
Lbot_589_590 bot589 bot590 {l}
Rtop_589_619 top589 top619 {r}
Ltop_589_619 top589 top619 {l}
Rbot_589_619 bot589 bot619 {r}
Lbot_589_619 bot589 bot619 {l}
C589 top589 bot589 {c}
Rtop_590_591 top590 top591 {r}
Ltop_590_591 top590 top591 {l}
Rbot_590_591 bot590 bot591 {r}
Lbot_590_591 bot590 bot591 {l}
Rtop_590_620 top590 top620 {r}
Ltop_590_620 top590 top620 {l}
Rbot_590_620 bot590 bot620 {r}
Lbot_590_620 bot590 bot620 {l}
C590 top590 bot590 {c}
Rtop_591_592 top591 top592 {r}
Ltop_591_592 top591 top592 {l}
Rbot_591_592 bot591 bot592 {r}
Lbot_591_592 bot591 bot592 {l}
Rtop_591_621 top591 top621 {r}
Ltop_591_621 top591 top621 {l}
Rbot_591_621 bot591 bot621 {r}
Lbot_591_621 bot591 bot621 {l}
C591 top591 bot591 {c}
Rtop_592_593 top592 top593 {r}
Ltop_592_593 top592 top593 {l}
Rbot_592_593 bot592 bot593 {r}
Lbot_592_593 bot592 bot593 {l}
Rtop_592_622 top592 top622 {r}
Ltop_592_622 top592 top622 {l}
Rbot_592_622 bot592 bot622 {r}
Lbot_592_622 bot592 bot622 {l}
C592 top592 bot592 {c}
Rtop_593_594 top593 top594 {r}
Ltop_593_594 top593 top594 {l}
Rbot_593_594 bot593 bot594 {r}
Lbot_593_594 bot593 bot594 {l}
Rtop_593_623 top593 top623 {r}
Ltop_593_623 top593 top623 {l}
Rbot_593_623 bot593 bot623 {r}
Lbot_593_623 bot593 bot623 {l}
C593 top593 bot593 {c}
Rtop_594_595 top594 top595 {r}
Ltop_594_595 top594 top595 {l}
Rbot_594_595 bot594 bot595 {r}
Lbot_594_595 bot594 bot595 {l}
Rtop_594_624 top594 top624 {r}
Ltop_594_624 top594 top624 {l}
Rbot_594_624 bot594 bot624 {r}
Lbot_594_624 bot594 bot624 {l}
C594 top594 bot594 {c}
Rtop_595_596 top595 top596 {r}
Ltop_595_596 top595 top596 {l}
Rbot_595_596 bot595 bot596 {r}
Lbot_595_596 bot595 bot596 {l}
Rtop_595_625 top595 top625 {r}
Ltop_595_625 top595 top625 {l}
Rbot_595_625 bot595 bot625 {r}
Lbot_595_625 bot595 bot625 {l}
C595 top595 bot595 {c}
Rtop_596_597 top596 top597 {r}
Ltop_596_597 top596 top597 {l}
Rbot_596_597 bot596 bot597 {r}
Lbot_596_597 bot596 bot597 {l}
Rtop_596_626 top596 top626 {r}
Ltop_596_626 top596 top626 {l}
Rbot_596_626 bot596 bot626 {r}
Lbot_596_626 bot596 bot626 {l}
C596 top596 bot596 {c}
Rtop_597_598 top597 top598 {r}
Ltop_597_598 top597 top598 {l}
Rbot_597_598 bot597 bot598 {r}
Lbot_597_598 bot597 bot598 {l}
Rtop_597_627 top597 top627 {r}
Ltop_597_627 top597 top627 {l}
Rbot_597_627 bot597 bot627 {r}
Lbot_597_627 bot597 bot627 {l}
C597 top597 bot597 {c}
Rtop_598_599 top598 top599 {r}
Ltop_598_599 top598 top599 {l}
Rbot_598_599 bot598 bot599 {r}
Lbot_598_599 bot598 bot599 {l}
Rtop_598_628 top598 top628 {r}
Ltop_598_628 top598 top628 {l}
Rbot_598_628 bot598 bot628 {r}
Lbot_598_628 bot598 bot628 {l}
C598 top598 bot598 {c}
Rtop_599_600 top599 top600 {r}
Ltop_599_600 top599 top600 {l}
Rbot_599_600 bot599 bot600 {r}
Lbot_599_600 bot599 bot600 {l}
Rtop_599_629 top599 top629 {r}
Ltop_599_629 top599 top629 {l}
Rbot_599_629 bot599 bot629 {r}
Lbot_599_629 bot599 bot629 {l}
C599 top599 bot599 {c}
Rtop_600_630 top600 top630 {r}
Ltop_600_630 top600 top630 {l}
Rbot_600_630 bot600 bot630 {r}
Lbot_600_630 bot600 bot630 {l}
C600 top600 bot600 {c}
Rtop_601_602 top601 top602 {r}
Ltop_601_602 top601 top602 {l}
Rbot_601_602 bot601 bot602 {r}
Lbot_601_602 bot601 bot602 {l}
Rtop_601_631 top601 top631 {r}
Ltop_601_631 top601 top631 {l}
Rbot_601_631 bot601 bot631 {r}
Lbot_601_631 bot601 bot631 {l}
C601 top601 bot601 {c}
Rtop_602_603 top602 top603 {r}
Ltop_602_603 top602 top603 {l}
Rbot_602_603 bot602 bot603 {r}
Lbot_602_603 bot602 bot603 {l}
Rtop_602_632 top602 top632 {r}
Ltop_602_632 top602 top632 {l}
Rbot_602_632 bot602 bot632 {r}
Lbot_602_632 bot602 bot632 {l}
C602 top602 bot602 {c}
Rtop_603_604 top603 top604 {r}
Ltop_603_604 top603 top604 {l}
Rbot_603_604 bot603 bot604 {r}
Lbot_603_604 bot603 bot604 {l}
Rtop_603_633 top603 top633 {r}
Ltop_603_633 top603 top633 {l}
Rbot_603_633 bot603 bot633 {r}
Lbot_603_633 bot603 bot633 {l}
C603 top603 bot603 {c}
Rtop_604_605 top604 top605 {r}
Ltop_604_605 top604 top605 {l}
Rbot_604_605 bot604 bot605 {r}
Lbot_604_605 bot604 bot605 {l}
Rtop_604_634 top604 top634 {r}
Ltop_604_634 top604 top634 {l}
Rbot_604_634 bot604 bot634 {r}
Lbot_604_634 bot604 bot634 {l}
C604 top604 bot604 {c}
Rtop_605_606 top605 top606 {r}
Ltop_605_606 top605 top606 {l}
Rbot_605_606 bot605 bot606 {r}
Lbot_605_606 bot605 bot606 {l}
Rtop_605_635 top605 top635 {r}
Ltop_605_635 top605 top635 {l}
Rbot_605_635 bot605 bot635 {r}
Lbot_605_635 bot605 bot635 {l}
C605 top605 bot605 {c}
Rtop_606_607 top606 top607 {r}
Ltop_606_607 top606 top607 {l}
Rbot_606_607 bot606 bot607 {r}
Lbot_606_607 bot606 bot607 {l}
Rtop_606_636 top606 top636 {r}
Ltop_606_636 top606 top636 {l}
Rbot_606_636 bot606 bot636 {r}
Lbot_606_636 bot606 bot636 {l}
C606 top606 bot606 {c}
Rtop_607_608 top607 top608 {r}
Ltop_607_608 top607 top608 {l}
Rbot_607_608 bot607 bot608 {r}
Lbot_607_608 bot607 bot608 {l}
Rtop_607_637 top607 top637 {r}
Ltop_607_637 top607 top637 {l}
Rbot_607_637 bot607 bot637 {r}
Lbot_607_637 bot607 bot637 {l}
C607 top607 bot607 {c}
Rtop_608_609 top608 top609 {r}
Ltop_608_609 top608 top609 {l}
Rbot_608_609 bot608 bot609 {r}
Lbot_608_609 bot608 bot609 {l}
Rtop_608_638 top608 top638 {r}
Ltop_608_638 top608 top638 {l}
Rbot_608_638 bot608 bot638 {r}
Lbot_608_638 bot608 bot638 {l}
C608 top608 bot608 {c}
Rtop_609_610 top609 top610 {r}
Ltop_609_610 top609 top610 {l}
Rbot_609_610 bot609 bot610 {r}
Lbot_609_610 bot609 bot610 {l}
Rtop_609_639 top609 top639 {r}
Ltop_609_639 top609 top639 {l}
Rbot_609_639 bot609 bot639 {r}
Lbot_609_639 bot609 bot639 {l}
C609 top609 bot609 {c}
Rtop_610_611 top610 top611 {r}
Ltop_610_611 top610 top611 {l}
Rbot_610_611 bot610 bot611 {r}
Lbot_610_611 bot610 bot611 {l}
Rtop_610_640 top610 top640 {r}
Ltop_610_640 top610 top640 {l}
Rbot_610_640 bot610 bot640 {r}
Lbot_610_640 bot610 bot640 {l}
C610 top610 bot610 {c}
Rtop_611_612 top611 top612 {r}
Ltop_611_612 top611 top612 {l}
Rbot_611_612 bot611 bot612 {r}
Lbot_611_612 bot611 bot612 {l}
Rtop_611_641 top611 top641 {r}
Ltop_611_641 top611 top641 {l}
Rbot_611_641 bot611 bot641 {r}
Lbot_611_641 bot611 bot641 {l}
C611 top611 bot611 {c}
Rtop_612_613 top612 top613 {r}
Ltop_612_613 top612 top613 {l}
Rbot_612_613 bot612 bot613 {r}
Lbot_612_613 bot612 bot613 {l}
Rtop_612_642 top612 top642 {r}
Ltop_612_642 top612 top642 {l}
Rbot_612_642 bot612 bot642 {r}
Lbot_612_642 bot612 bot642 {l}
C612 top612 bot612 {c}
Rtop_613_614 top613 top614 {r}
Ltop_613_614 top613 top614 {l}
Rbot_613_614 bot613 bot614 {r}
Lbot_613_614 bot613 bot614 {l}
Rtop_613_643 top613 top643 {r}
Ltop_613_643 top613 top643 {l}
Rbot_613_643 bot613 bot643 {r}
Lbot_613_643 bot613 bot643 {l}
C613 top613 bot613 {c}
Rtop_614_615 top614 top615 {r}
Ltop_614_615 top614 top615 {l}
Rbot_614_615 bot614 bot615 {r}
Lbot_614_615 bot614 bot615 {l}
Rtop_614_644 top614 top644 {r}
Ltop_614_644 top614 top644 {l}
Rbot_614_644 bot614 bot644 {r}
Lbot_614_644 bot614 bot644 {l}
C614 top614 bot614 {c}
Rtop_615_616 top615 top616 {r}
Ltop_615_616 top615 top616 {l}
Rbot_615_616 bot615 bot616 {r}
Lbot_615_616 bot615 bot616 {l}
Rtop_615_645 top615 top645 {r}
Ltop_615_645 top615 top645 {l}
Rbot_615_645 bot615 bot645 {r}
Lbot_615_645 bot615 bot645 {l}
C615 top615 bot615 {c}
Rtop_616_617 top616 top617 {r}
Ltop_616_617 top616 top617 {l}
Rbot_616_617 bot616 bot617 {r}
Lbot_616_617 bot616 bot617 {l}
Rtop_616_646 top616 top646 {r}
Ltop_616_646 top616 top646 {l}
Rbot_616_646 bot616 bot646 {r}
Lbot_616_646 bot616 bot646 {l}
C616 top616 bot616 {c}
Rtop_617_618 top617 top618 {r}
Ltop_617_618 top617 top618 {l}
Rbot_617_618 bot617 bot618 {r}
Lbot_617_618 bot617 bot618 {l}
Rtop_617_647 top617 top647 {r}
Ltop_617_647 top617 top647 {l}
Rbot_617_647 bot617 bot647 {r}
Lbot_617_647 bot617 bot647 {l}
C617 top617 bot617 {c}
Rtop_618_619 top618 top619 {r}
Ltop_618_619 top618 top619 {l}
Rbot_618_619 bot618 bot619 {r}
Lbot_618_619 bot618 bot619 {l}
Rtop_618_648 top618 top648 {r}
Ltop_618_648 top618 top648 {l}
Rbot_618_648 bot618 bot648 {r}
Lbot_618_648 bot618 bot648 {l}
C618 top618 bot618 {c}
Rtop_619_620 top619 top620 {r}
Ltop_619_620 top619 top620 {l}
Rbot_619_620 bot619 bot620 {r}
Lbot_619_620 bot619 bot620 {l}
Rtop_619_649 top619 top649 {r}
Ltop_619_649 top619 top649 {l}
Rbot_619_649 bot619 bot649 {r}
Lbot_619_649 bot619 bot649 {l}
C619 top619 bot619 {c}
Rtop_620_621 top620 top621 {r}
Ltop_620_621 top620 top621 {l}
Rbot_620_621 bot620 bot621 {r}
Lbot_620_621 bot620 bot621 {l}
Rtop_620_650 top620 top650 {r}
Ltop_620_650 top620 top650 {l}
Rbot_620_650 bot620 bot650 {r}
Lbot_620_650 bot620 bot650 {l}
C620 top620 bot620 {c}
Rtop_621_622 top621 top622 {r}
Ltop_621_622 top621 top622 {l}
Rbot_621_622 bot621 bot622 {r}
Lbot_621_622 bot621 bot622 {l}
Rtop_621_651 top621 top651 {r}
Ltop_621_651 top621 top651 {l}
Rbot_621_651 bot621 bot651 {r}
Lbot_621_651 bot621 bot651 {l}
C621 top621 bot621 {c}
Rtop_622_623 top622 top623 {r}
Ltop_622_623 top622 top623 {l}
Rbot_622_623 bot622 bot623 {r}
Lbot_622_623 bot622 bot623 {l}
Rtop_622_652 top622 top652 {r}
Ltop_622_652 top622 top652 {l}
Rbot_622_652 bot622 bot652 {r}
Lbot_622_652 bot622 bot652 {l}
C622 top622 bot622 {c}
Rtop_623_624 top623 top624 {r}
Ltop_623_624 top623 top624 {l}
Rbot_623_624 bot623 bot624 {r}
Lbot_623_624 bot623 bot624 {l}
Rtop_623_653 top623 top653 {r}
Ltop_623_653 top623 top653 {l}
Rbot_623_653 bot623 bot653 {r}
Lbot_623_653 bot623 bot653 {l}
C623 top623 bot623 {c}
Rtop_624_625 top624 top625 {r}
Ltop_624_625 top624 top625 {l}
Rbot_624_625 bot624 bot625 {r}
Lbot_624_625 bot624 bot625 {l}
Rtop_624_654 top624 top654 {r}
Ltop_624_654 top624 top654 {l}
Rbot_624_654 bot624 bot654 {r}
Lbot_624_654 bot624 bot654 {l}
C624 top624 bot624 {c}
Rtop_625_626 top625 top626 {r}
Ltop_625_626 top625 top626 {l}
Rbot_625_626 bot625 bot626 {r}
Lbot_625_626 bot625 bot626 {l}
Rtop_625_655 top625 top655 {r}
Ltop_625_655 top625 top655 {l}
Rbot_625_655 bot625 bot655 {r}
Lbot_625_655 bot625 bot655 {l}
C625 top625 bot625 {c}
Rtop_626_627 top626 top627 {r}
Ltop_626_627 top626 top627 {l}
Rbot_626_627 bot626 bot627 {r}
Lbot_626_627 bot626 bot627 {l}
Rtop_626_656 top626 top656 {r}
Ltop_626_656 top626 top656 {l}
Rbot_626_656 bot626 bot656 {r}
Lbot_626_656 bot626 bot656 {l}
C626 top626 bot626 {c}
Rtop_627_628 top627 top628 {r}
Ltop_627_628 top627 top628 {l}
Rbot_627_628 bot627 bot628 {r}
Lbot_627_628 bot627 bot628 {l}
Rtop_627_657 top627 top657 {r}
Ltop_627_657 top627 top657 {l}
Rbot_627_657 bot627 bot657 {r}
Lbot_627_657 bot627 bot657 {l}
C627 top627 bot627 {c}
Rtop_628_629 top628 top629 {r}
Ltop_628_629 top628 top629 {l}
Rbot_628_629 bot628 bot629 {r}
Lbot_628_629 bot628 bot629 {l}
Rtop_628_658 top628 top658 {r}
Ltop_628_658 top628 top658 {l}
Rbot_628_658 bot628 bot658 {r}
Lbot_628_658 bot628 bot658 {l}
C628 top628 bot628 {c}
Rtop_629_630 top629 top630 {r}
Ltop_629_630 top629 top630 {l}
Rbot_629_630 bot629 bot630 {r}
Lbot_629_630 bot629 bot630 {l}
Rtop_629_659 top629 top659 {r}
Ltop_629_659 top629 top659 {l}
Rbot_629_659 bot629 bot659 {r}
Lbot_629_659 bot629 bot659 {l}
C629 top629 bot629 {c}
Rtop_630_660 top630 top660 {r}
Ltop_630_660 top630 top660 {l}
Rbot_630_660 bot630 bot660 {r}
Lbot_630_660 bot630 bot660 {l}
C630 top630 bot630 {c}
Rtop_631_632 top631 top632 {r}
Ltop_631_632 top631 top632 {l}
Rbot_631_632 bot631 bot632 {r}
Lbot_631_632 bot631 bot632 {l}
Rtop_631_661 top631 top661 {r}
Ltop_631_661 top631 top661 {l}
Rbot_631_661 bot631 bot661 {r}
Lbot_631_661 bot631 bot661 {l}
C631 top631 bot631 {c}
Rtop_632_633 top632 top633 {r}
Ltop_632_633 top632 top633 {l}
Rbot_632_633 bot632 bot633 {r}
Lbot_632_633 bot632 bot633 {l}
Rtop_632_662 top632 top662 {r}
Ltop_632_662 top632 top662 {l}
Rbot_632_662 bot632 bot662 {r}
Lbot_632_662 bot632 bot662 {l}
C632 top632 bot632 {c}
Rtop_633_634 top633 top634 {r}
Ltop_633_634 top633 top634 {l}
Rbot_633_634 bot633 bot634 {r}
Lbot_633_634 bot633 bot634 {l}
Rtop_633_663 top633 top663 {r}
Ltop_633_663 top633 top663 {l}
Rbot_633_663 bot633 bot663 {r}
Lbot_633_663 bot633 bot663 {l}
C633 top633 bot633 {c}
Rtop_634_635 top634 top635 {r}
Ltop_634_635 top634 top635 {l}
Rbot_634_635 bot634 bot635 {r}
Lbot_634_635 bot634 bot635 {l}
Rtop_634_664 top634 top664 {r}
Ltop_634_664 top634 top664 {l}
Rbot_634_664 bot634 bot664 {r}
Lbot_634_664 bot634 bot664 {l}
C634 top634 bot634 {c}
Rtop_635_636 top635 top636 {r}
Ltop_635_636 top635 top636 {l}
Rbot_635_636 bot635 bot636 {r}
Lbot_635_636 bot635 bot636 {l}
Rtop_635_665 top635 top665 {r}
Ltop_635_665 top635 top665 {l}
Rbot_635_665 bot635 bot665 {r}
Lbot_635_665 bot635 bot665 {l}
C635 top635 bot635 {c}
Rtop_636_637 top636 top637 {r}
Ltop_636_637 top636 top637 {l}
Rbot_636_637 bot636 bot637 {r}
Lbot_636_637 bot636 bot637 {l}
Rtop_636_666 top636 top666 {r}
Ltop_636_666 top636 top666 {l}
Rbot_636_666 bot636 bot666 {r}
Lbot_636_666 bot636 bot666 {l}
C636 top636 bot636 {c}
Rtop_637_638 top637 top638 {r}
Ltop_637_638 top637 top638 {l}
Rbot_637_638 bot637 bot638 {r}
Lbot_637_638 bot637 bot638 {l}
Rtop_637_667 top637 top667 {r}
Ltop_637_667 top637 top667 {l}
Rbot_637_667 bot637 bot667 {r}
Lbot_637_667 bot637 bot667 {l}
C637 top637 bot637 {c}
Rtop_638_639 top638 top639 {r}
Ltop_638_639 top638 top639 {l}
Rbot_638_639 bot638 bot639 {r}
Lbot_638_639 bot638 bot639 {l}
Rtop_638_668 top638 top668 {r}
Ltop_638_668 top638 top668 {l}
Rbot_638_668 bot638 bot668 {r}
Lbot_638_668 bot638 bot668 {l}
C638 top638 bot638 {c}
Rtop_639_640 top639 top640 {r}
Ltop_639_640 top639 top640 {l}
Rbot_639_640 bot639 bot640 {r}
Lbot_639_640 bot639 bot640 {l}
Rtop_639_669 top639 top669 {r}
Ltop_639_669 top639 top669 {l}
Rbot_639_669 bot639 bot669 {r}
Lbot_639_669 bot639 bot669 {l}
C639 top639 bot639 {c}
Rtop_640_641 top640 top641 {r}
Ltop_640_641 top640 top641 {l}
Rbot_640_641 bot640 bot641 {r}
Lbot_640_641 bot640 bot641 {l}
Rtop_640_670 top640 top670 {r}
Ltop_640_670 top640 top670 {l}
Rbot_640_670 bot640 bot670 {r}
Lbot_640_670 bot640 bot670 {l}
C640 top640 bot640 {c}
Rtop_641_642 top641 top642 {r}
Ltop_641_642 top641 top642 {l}
Rbot_641_642 bot641 bot642 {r}
Lbot_641_642 bot641 bot642 {l}
Rtop_641_671 top641 top671 {r}
Ltop_641_671 top641 top671 {l}
Rbot_641_671 bot641 bot671 {r}
Lbot_641_671 bot641 bot671 {l}
C641 top641 bot641 {c}
Rtop_642_643 top642 top643 {r}
Ltop_642_643 top642 top643 {l}
Rbot_642_643 bot642 bot643 {r}
Lbot_642_643 bot642 bot643 {l}
Rtop_642_672 top642 top672 {r}
Ltop_642_672 top642 top672 {l}
Rbot_642_672 bot642 bot672 {r}
Lbot_642_672 bot642 bot672 {l}
C642 top642 bot642 {c}
Rtop_643_644 top643 top644 {r}
Ltop_643_644 top643 top644 {l}
Rbot_643_644 bot643 bot644 {r}
Lbot_643_644 bot643 bot644 {l}
Rtop_643_673 top643 top673 {r}
Ltop_643_673 top643 top673 {l}
Rbot_643_673 bot643 bot673 {r}
Lbot_643_673 bot643 bot673 {l}
C643 top643 bot643 {c}
Rtop_644_645 top644 top645 {r}
Ltop_644_645 top644 top645 {l}
Rbot_644_645 bot644 bot645 {r}
Lbot_644_645 bot644 bot645 {l}
Rtop_644_674 top644 top674 {r}
Ltop_644_674 top644 top674 {l}
Rbot_644_674 bot644 bot674 {r}
Lbot_644_674 bot644 bot674 {l}
C644 top644 bot644 {c}
Rtop_645_646 top645 top646 {r}
Ltop_645_646 top645 top646 {l}
Rbot_645_646 bot645 bot646 {r}
Lbot_645_646 bot645 bot646 {l}
Rtop_645_675 top645 top675 {r}
Ltop_645_675 top645 top675 {l}
Rbot_645_675 bot645 bot675 {r}
Lbot_645_675 bot645 bot675 {l}
C645 top645 bot645 {c}
Rtop_646_647 top646 top647 {r}
Ltop_646_647 top646 top647 {l}
Rbot_646_647 bot646 bot647 {r}
Lbot_646_647 bot646 bot647 {l}
Rtop_646_676 top646 top676 {r}
Ltop_646_676 top646 top676 {l}
Rbot_646_676 bot646 bot676 {r}
Lbot_646_676 bot646 bot676 {l}
C646 top646 bot646 {c}
Rtop_647_648 top647 top648 {r}
Ltop_647_648 top647 top648 {l}
Rbot_647_648 bot647 bot648 {r}
Lbot_647_648 bot647 bot648 {l}
Rtop_647_677 top647 top677 {r}
Ltop_647_677 top647 top677 {l}
Rbot_647_677 bot647 bot677 {r}
Lbot_647_677 bot647 bot677 {l}
C647 top647 bot647 {c}
Rtop_648_649 top648 top649 {r}
Ltop_648_649 top648 top649 {l}
Rbot_648_649 bot648 bot649 {r}
Lbot_648_649 bot648 bot649 {l}
Rtop_648_678 top648 top678 {r}
Ltop_648_678 top648 top678 {l}
Rbot_648_678 bot648 bot678 {r}
Lbot_648_678 bot648 bot678 {l}
C648 top648 bot648 {c}
Rtop_649_650 top649 top650 {r}
Ltop_649_650 top649 top650 {l}
Rbot_649_650 bot649 bot650 {r}
Lbot_649_650 bot649 bot650 {l}
Rtop_649_679 top649 top679 {r}
Ltop_649_679 top649 top679 {l}
Rbot_649_679 bot649 bot679 {r}
Lbot_649_679 bot649 bot679 {l}
C649 top649 bot649 {c}
Rtop_650_651 top650 top651 {r}
Ltop_650_651 top650 top651 {l}
Rbot_650_651 bot650 bot651 {r}
Lbot_650_651 bot650 bot651 {l}
Rtop_650_680 top650 top680 {r}
Ltop_650_680 top650 top680 {l}
Rbot_650_680 bot650 bot680 {r}
Lbot_650_680 bot650 bot680 {l}
C650 top650 bot650 {c}
Rtop_651_652 top651 top652 {r}
Ltop_651_652 top651 top652 {l}
Rbot_651_652 bot651 bot652 {r}
Lbot_651_652 bot651 bot652 {l}
Rtop_651_681 top651 top681 {r}
Ltop_651_681 top651 top681 {l}
Rbot_651_681 bot651 bot681 {r}
Lbot_651_681 bot651 bot681 {l}
C651 top651 bot651 {c}
Rtop_652_653 top652 top653 {r}
Ltop_652_653 top652 top653 {l}
Rbot_652_653 bot652 bot653 {r}
Lbot_652_653 bot652 bot653 {l}
Rtop_652_682 top652 top682 {r}
Ltop_652_682 top652 top682 {l}
Rbot_652_682 bot652 bot682 {r}
Lbot_652_682 bot652 bot682 {l}
C652 top652 bot652 {c}
Rtop_653_654 top653 top654 {r}
Ltop_653_654 top653 top654 {l}
Rbot_653_654 bot653 bot654 {r}
Lbot_653_654 bot653 bot654 {l}
Rtop_653_683 top653 top683 {r}
Ltop_653_683 top653 top683 {l}
Rbot_653_683 bot653 bot683 {r}
Lbot_653_683 bot653 bot683 {l}
C653 top653 bot653 {c}
Rtop_654_655 top654 top655 {r}
Ltop_654_655 top654 top655 {l}
Rbot_654_655 bot654 bot655 {r}
Lbot_654_655 bot654 bot655 {l}
Rtop_654_684 top654 top684 {r}
Ltop_654_684 top654 top684 {l}
Rbot_654_684 bot654 bot684 {r}
Lbot_654_684 bot654 bot684 {l}
C654 top654 bot654 {c}
Rtop_655_656 top655 top656 {r}
Ltop_655_656 top655 top656 {l}
Rbot_655_656 bot655 bot656 {r}
Lbot_655_656 bot655 bot656 {l}
Rtop_655_685 top655 top685 {r}
Ltop_655_685 top655 top685 {l}
Rbot_655_685 bot655 bot685 {r}
Lbot_655_685 bot655 bot685 {l}
C655 top655 bot655 {c}
Rtop_656_657 top656 top657 {r}
Ltop_656_657 top656 top657 {l}
Rbot_656_657 bot656 bot657 {r}
Lbot_656_657 bot656 bot657 {l}
Rtop_656_686 top656 top686 {r}
Ltop_656_686 top656 top686 {l}
Rbot_656_686 bot656 bot686 {r}
Lbot_656_686 bot656 bot686 {l}
C656 top656 bot656 {c}
Rtop_657_658 top657 top658 {r}
Ltop_657_658 top657 top658 {l}
Rbot_657_658 bot657 bot658 {r}
Lbot_657_658 bot657 bot658 {l}
Rtop_657_687 top657 top687 {r}
Ltop_657_687 top657 top687 {l}
Rbot_657_687 bot657 bot687 {r}
Lbot_657_687 bot657 bot687 {l}
C657 top657 bot657 {c}
Rtop_658_659 top658 top659 {r}
Ltop_658_659 top658 top659 {l}
Rbot_658_659 bot658 bot659 {r}
Lbot_658_659 bot658 bot659 {l}
Rtop_658_688 top658 top688 {r}
Ltop_658_688 top658 top688 {l}
Rbot_658_688 bot658 bot688 {r}
Lbot_658_688 bot658 bot688 {l}
C658 top658 bot658 {c}
Rtop_659_660 top659 top660 {r}
Ltop_659_660 top659 top660 {l}
Rbot_659_660 bot659 bot660 {r}
Lbot_659_660 bot659 bot660 {l}
Rtop_659_689 top659 top689 {r}
Ltop_659_689 top659 top689 {l}
Rbot_659_689 bot659 bot689 {r}
Lbot_659_689 bot659 bot689 {l}
C659 top659 bot659 {c}
Rtop_660_690 top660 top690 {r}
Ltop_660_690 top660 top690 {l}
Rbot_660_690 bot660 bot690 {r}
Lbot_660_690 bot660 bot690 {l}
C660 top660 bot660 {c}
Rtop_661_662 top661 top662 {r}
Ltop_661_662 top661 top662 {l}
Rbot_661_662 bot661 bot662 {r}
Lbot_661_662 bot661 bot662 {l}
Rtop_661_691 top661 top691 {r}
Ltop_661_691 top661 top691 {l}
Rbot_661_691 bot661 bot691 {r}
Lbot_661_691 bot661 bot691 {l}
C661 top661 bot661 {c}
Rtop_662_663 top662 top663 {r}
Ltop_662_663 top662 top663 {l}
Rbot_662_663 bot662 bot663 {r}
Lbot_662_663 bot662 bot663 {l}
Rtop_662_692 top662 top692 {r}
Ltop_662_692 top662 top692 {l}
Rbot_662_692 bot662 bot692 {r}
Lbot_662_692 bot662 bot692 {l}
C662 top662 bot662 {c}
Rtop_663_664 top663 top664 {r}
Ltop_663_664 top663 top664 {l}
Rbot_663_664 bot663 bot664 {r}
Lbot_663_664 bot663 bot664 {l}
Rtop_663_693 top663 top693 {r}
Ltop_663_693 top663 top693 {l}
Rbot_663_693 bot663 bot693 {r}
Lbot_663_693 bot663 bot693 {l}
C663 top663 bot663 {c}
Rtop_664_665 top664 top665 {r}
Ltop_664_665 top664 top665 {l}
Rbot_664_665 bot664 bot665 {r}
Lbot_664_665 bot664 bot665 {l}
Rtop_664_694 top664 top694 {r}
Ltop_664_694 top664 top694 {l}
Rbot_664_694 bot664 bot694 {r}
Lbot_664_694 bot664 bot694 {l}
C664 top664 bot664 {c}
Rtop_665_666 top665 top666 {r}
Ltop_665_666 top665 top666 {l}
Rbot_665_666 bot665 bot666 {r}
Lbot_665_666 bot665 bot666 {l}
Rtop_665_695 top665 top695 {r}
Ltop_665_695 top665 top695 {l}
Rbot_665_695 bot665 bot695 {r}
Lbot_665_695 bot665 bot695 {l}
C665 top665 bot665 {c}
Rtop_666_667 top666 top667 {r}
Ltop_666_667 top666 top667 {l}
Rbot_666_667 bot666 bot667 {r}
Lbot_666_667 bot666 bot667 {l}
Rtop_666_696 top666 top696 {r}
Ltop_666_696 top666 top696 {l}
Rbot_666_696 bot666 bot696 {r}
Lbot_666_696 bot666 bot696 {l}
C666 top666 bot666 {c}
Rtop_667_668 top667 top668 {r}
Ltop_667_668 top667 top668 {l}
Rbot_667_668 bot667 bot668 {r}
Lbot_667_668 bot667 bot668 {l}
Rtop_667_697 top667 top697 {r}
Ltop_667_697 top667 top697 {l}
Rbot_667_697 bot667 bot697 {r}
Lbot_667_697 bot667 bot697 {l}
C667 top667 bot667 {c}
Rtop_668_669 top668 top669 {r}
Ltop_668_669 top668 top669 {l}
Rbot_668_669 bot668 bot669 {r}
Lbot_668_669 bot668 bot669 {l}
Rtop_668_698 top668 top698 {r}
Ltop_668_698 top668 top698 {l}
Rbot_668_698 bot668 bot698 {r}
Lbot_668_698 bot668 bot698 {l}
C668 top668 bot668 {c}
Rtop_669_670 top669 top670 {r}
Ltop_669_670 top669 top670 {l}
Rbot_669_670 bot669 bot670 {r}
Lbot_669_670 bot669 bot670 {l}
Rtop_669_699 top669 top699 {r}
Ltop_669_699 top669 top699 {l}
Rbot_669_699 bot669 bot699 {r}
Lbot_669_699 bot669 bot699 {l}
C669 top669 bot669 {c}
Rtop_670_671 top670 top671 {r}
Ltop_670_671 top670 top671 {l}
Rbot_670_671 bot670 bot671 {r}
Lbot_670_671 bot670 bot671 {l}
Rtop_670_700 top670 top700 {r}
Ltop_670_700 top670 top700 {l}
Rbot_670_700 bot670 bot700 {r}
Lbot_670_700 bot670 bot700 {l}
C670 top670 bot670 {c}
Rtop_671_672 top671 top672 {r}
Ltop_671_672 top671 top672 {l}
Rbot_671_672 bot671 bot672 {r}
Lbot_671_672 bot671 bot672 {l}
Rtop_671_701 top671 top701 {r}
Ltop_671_701 top671 top701 {l}
Rbot_671_701 bot671 bot701 {r}
Lbot_671_701 bot671 bot701 {l}
C671 top671 bot671 {c}
Rtop_672_673 top672 top673 {r}
Ltop_672_673 top672 top673 {l}
Rbot_672_673 bot672 bot673 {r}
Lbot_672_673 bot672 bot673 {l}
Rtop_672_702 top672 top702 {r}
Ltop_672_702 top672 top702 {l}
Rbot_672_702 bot672 bot702 {r}
Lbot_672_702 bot672 bot702 {l}
C672 top672 bot672 {c}
Rtop_673_674 top673 top674 {r}
Ltop_673_674 top673 top674 {l}
Rbot_673_674 bot673 bot674 {r}
Lbot_673_674 bot673 bot674 {l}
Rtop_673_703 top673 top703 {r}
Ltop_673_703 top673 top703 {l}
Rbot_673_703 bot673 bot703 {r}
Lbot_673_703 bot673 bot703 {l}
C673 top673 bot673 {c}
Rtop_674_675 top674 top675 {r}
Ltop_674_675 top674 top675 {l}
Rbot_674_675 bot674 bot675 {r}
Lbot_674_675 bot674 bot675 {l}
Rtop_674_704 top674 top704 {r}
Ltop_674_704 top674 top704 {l}
Rbot_674_704 bot674 bot704 {r}
Lbot_674_704 bot674 bot704 {l}
C674 top674 bot674 {c}
Rtop_675_676 top675 top676 {r}
Ltop_675_676 top675 top676 {l}
Rbot_675_676 bot675 bot676 {r}
Lbot_675_676 bot675 bot676 {l}
Rtop_675_705 top675 top705 {r}
Ltop_675_705 top675 top705 {l}
Rbot_675_705 bot675 bot705 {r}
Lbot_675_705 bot675 bot705 {l}
C675 top675 bot675 {c}
Rtop_676_677 top676 top677 {r}
Ltop_676_677 top676 top677 {l}
Rbot_676_677 bot676 bot677 {r}
Lbot_676_677 bot676 bot677 {l}
Rtop_676_706 top676 top706 {r}
Ltop_676_706 top676 top706 {l}
Rbot_676_706 bot676 bot706 {r}
Lbot_676_706 bot676 bot706 {l}
C676 top676 bot676 {c}
Rtop_677_678 top677 top678 {r}
Ltop_677_678 top677 top678 {l}
Rbot_677_678 bot677 bot678 {r}
Lbot_677_678 bot677 bot678 {l}
Rtop_677_707 top677 top707 {r}
Ltop_677_707 top677 top707 {l}
Rbot_677_707 bot677 bot707 {r}
Lbot_677_707 bot677 bot707 {l}
C677 top677 bot677 {c}
Rtop_678_679 top678 top679 {r}
Ltop_678_679 top678 top679 {l}
Rbot_678_679 bot678 bot679 {r}
Lbot_678_679 bot678 bot679 {l}
Rtop_678_708 top678 top708 {r}
Ltop_678_708 top678 top708 {l}
Rbot_678_708 bot678 bot708 {r}
Lbot_678_708 bot678 bot708 {l}
C678 top678 bot678 {c}
Rtop_679_680 top679 top680 {r}
Ltop_679_680 top679 top680 {l}
Rbot_679_680 bot679 bot680 {r}
Lbot_679_680 bot679 bot680 {l}
Rtop_679_709 top679 top709 {r}
Ltop_679_709 top679 top709 {l}
Rbot_679_709 bot679 bot709 {r}
Lbot_679_709 bot679 bot709 {l}
C679 top679 bot679 {c}
Rtop_680_681 top680 top681 {r}
Ltop_680_681 top680 top681 {l}
Rbot_680_681 bot680 bot681 {r}
Lbot_680_681 bot680 bot681 {l}
Rtop_680_710 top680 top710 {r}
Ltop_680_710 top680 top710 {l}
Rbot_680_710 bot680 bot710 {r}
Lbot_680_710 bot680 bot710 {l}
C680 top680 bot680 {c}
Rtop_681_682 top681 top682 {r}
Ltop_681_682 top681 top682 {l}
Rbot_681_682 bot681 bot682 {r}
Lbot_681_682 bot681 bot682 {l}
Rtop_681_711 top681 top711 {r}
Ltop_681_711 top681 top711 {l}
Rbot_681_711 bot681 bot711 {r}
Lbot_681_711 bot681 bot711 {l}
C681 top681 bot681 {c}
Rtop_682_683 top682 top683 {r}
Ltop_682_683 top682 top683 {l}
Rbot_682_683 bot682 bot683 {r}
Lbot_682_683 bot682 bot683 {l}
Rtop_682_712 top682 top712 {r}
Ltop_682_712 top682 top712 {l}
Rbot_682_712 bot682 bot712 {r}
Lbot_682_712 bot682 bot712 {l}
C682 top682 bot682 {c}
Rtop_683_684 top683 top684 {r}
Ltop_683_684 top683 top684 {l}
Rbot_683_684 bot683 bot684 {r}
Lbot_683_684 bot683 bot684 {l}
Rtop_683_713 top683 top713 {r}
Ltop_683_713 top683 top713 {l}
Rbot_683_713 bot683 bot713 {r}
Lbot_683_713 bot683 bot713 {l}
C683 top683 bot683 {c}
Rtop_684_685 top684 top685 {r}
Ltop_684_685 top684 top685 {l}
Rbot_684_685 bot684 bot685 {r}
Lbot_684_685 bot684 bot685 {l}
Rtop_684_714 top684 top714 {r}
Ltop_684_714 top684 top714 {l}
Rbot_684_714 bot684 bot714 {r}
Lbot_684_714 bot684 bot714 {l}
C684 top684 bot684 {c}
Rtop_685_686 top685 top686 {r}
Ltop_685_686 top685 top686 {l}
Rbot_685_686 bot685 bot686 {r}
Lbot_685_686 bot685 bot686 {l}
Rtop_685_715 top685 top715 {r}
Ltop_685_715 top685 top715 {l}
Rbot_685_715 bot685 bot715 {r}
Lbot_685_715 bot685 bot715 {l}
C685 top685 bot685 {c}
Rtop_686_687 top686 top687 {r}
Ltop_686_687 top686 top687 {l}
Rbot_686_687 bot686 bot687 {r}
Lbot_686_687 bot686 bot687 {l}
Rtop_686_716 top686 top716 {r}
Ltop_686_716 top686 top716 {l}
Rbot_686_716 bot686 bot716 {r}
Lbot_686_716 bot686 bot716 {l}
C686 top686 bot686 {c}
Rtop_687_688 top687 top688 {r}
Ltop_687_688 top687 top688 {l}
Rbot_687_688 bot687 bot688 {r}
Lbot_687_688 bot687 bot688 {l}
Rtop_687_717 top687 top717 {r}
Ltop_687_717 top687 top717 {l}
Rbot_687_717 bot687 bot717 {r}
Lbot_687_717 bot687 bot717 {l}
C687 top687 bot687 {c}
Rtop_688_689 top688 top689 {r}
Ltop_688_689 top688 top689 {l}
Rbot_688_689 bot688 bot689 {r}
Lbot_688_689 bot688 bot689 {l}
Rtop_688_718 top688 top718 {r}
Ltop_688_718 top688 top718 {l}
Rbot_688_718 bot688 bot718 {r}
Lbot_688_718 bot688 bot718 {l}
C688 top688 bot688 {c}
Rtop_689_690 top689 top690 {r}
Ltop_689_690 top689 top690 {l}
Rbot_689_690 bot689 bot690 {r}
Lbot_689_690 bot689 bot690 {l}
Rtop_689_719 top689 top719 {r}
Ltop_689_719 top689 top719 {l}
Rbot_689_719 bot689 bot719 {r}
Lbot_689_719 bot689 bot719 {l}
C689 top689 bot689 {c}
Rtop_690_720 top690 top720 {r}
Ltop_690_720 top690 top720 {l}
Rbot_690_720 bot690 bot720 {r}
Lbot_690_720 bot690 bot720 {l}
C690 top690 bot690 {c}
Rtop_691_692 top691 top692 {r}
Ltop_691_692 top691 top692 {l}
Rbot_691_692 bot691 bot692 {r}
Lbot_691_692 bot691 bot692 {l}
Rtop_691_721 top691 top721 {r}
Ltop_691_721 top691 top721 {l}
Rbot_691_721 bot691 bot721 {r}
Lbot_691_721 bot691 bot721 {l}
C691 top691 bot691 {c}
Rtop_692_693 top692 top693 {r}
Ltop_692_693 top692 top693 {l}
Rbot_692_693 bot692 bot693 {r}
Lbot_692_693 bot692 bot693 {l}
Rtop_692_722 top692 top722 {r}
Ltop_692_722 top692 top722 {l}
Rbot_692_722 bot692 bot722 {r}
Lbot_692_722 bot692 bot722 {l}
C692 top692 bot692 {c}
Rtop_693_694 top693 top694 {r}
Ltop_693_694 top693 top694 {l}
Rbot_693_694 bot693 bot694 {r}
Lbot_693_694 bot693 bot694 {l}
Rtop_693_723 top693 top723 {r}
Ltop_693_723 top693 top723 {l}
Rbot_693_723 bot693 bot723 {r}
Lbot_693_723 bot693 bot723 {l}
C693 top693 bot693 {c}
Rtop_694_695 top694 top695 {r}
Ltop_694_695 top694 top695 {l}
Rbot_694_695 bot694 bot695 {r}
Lbot_694_695 bot694 bot695 {l}
Rtop_694_724 top694 top724 {r}
Ltop_694_724 top694 top724 {l}
Rbot_694_724 bot694 bot724 {r}
Lbot_694_724 bot694 bot724 {l}
C694 top694 bot694 {c}
Rtop_695_696 top695 top696 {r}
Ltop_695_696 top695 top696 {l}
Rbot_695_696 bot695 bot696 {r}
Lbot_695_696 bot695 bot696 {l}
Rtop_695_725 top695 top725 {r}
Ltop_695_725 top695 top725 {l}
Rbot_695_725 bot695 bot725 {r}
Lbot_695_725 bot695 bot725 {l}
C695 top695 bot695 {c}
Rtop_696_697 top696 top697 {r}
Ltop_696_697 top696 top697 {l}
Rbot_696_697 bot696 bot697 {r}
Lbot_696_697 bot696 bot697 {l}
Rtop_696_726 top696 top726 {r}
Ltop_696_726 top696 top726 {l}
Rbot_696_726 bot696 bot726 {r}
Lbot_696_726 bot696 bot726 {l}
C696 top696 bot696 {c}
Rtop_697_698 top697 top698 {r}
Ltop_697_698 top697 top698 {l}
Rbot_697_698 bot697 bot698 {r}
Lbot_697_698 bot697 bot698 {l}
Rtop_697_727 top697 top727 {r}
Ltop_697_727 top697 top727 {l}
Rbot_697_727 bot697 bot727 {r}
Lbot_697_727 bot697 bot727 {l}
C697 top697 bot697 {c}
Rtop_698_699 top698 top699 {r}
Ltop_698_699 top698 top699 {l}
Rbot_698_699 bot698 bot699 {r}
Lbot_698_699 bot698 bot699 {l}
Rtop_698_728 top698 top728 {r}
Ltop_698_728 top698 top728 {l}
Rbot_698_728 bot698 bot728 {r}
Lbot_698_728 bot698 bot728 {l}
C698 top698 bot698 {c}
Rtop_699_700 top699 top700 {r}
Ltop_699_700 top699 top700 {l}
Rbot_699_700 bot699 bot700 {r}
Lbot_699_700 bot699 bot700 {l}
Rtop_699_729 top699 top729 {r}
Ltop_699_729 top699 top729 {l}
Rbot_699_729 bot699 bot729 {r}
Lbot_699_729 bot699 bot729 {l}
C699 top699 bot699 {c}
Rtop_700_701 top700 top701 {r}
Ltop_700_701 top700 top701 {l}
Rbot_700_701 bot700 bot701 {r}
Lbot_700_701 bot700 bot701 {l}
Rtop_700_730 top700 top730 {r}
Ltop_700_730 top700 top730 {l}
Rbot_700_730 bot700 bot730 {r}
Lbot_700_730 bot700 bot730 {l}
C700 top700 bot700 {c}
Rtop_701_702 top701 top702 {r}
Ltop_701_702 top701 top702 {l}
Rbot_701_702 bot701 bot702 {r}
Lbot_701_702 bot701 bot702 {l}
Rtop_701_731 top701 top731 {r}
Ltop_701_731 top701 top731 {l}
Rbot_701_731 bot701 bot731 {r}
Lbot_701_731 bot701 bot731 {l}
C701 top701 bot701 {c}
Rtop_702_703 top702 top703 {r}
Ltop_702_703 top702 top703 {l}
Rbot_702_703 bot702 bot703 {r}
Lbot_702_703 bot702 bot703 {l}
Rtop_702_732 top702 top732 {r}
Ltop_702_732 top702 top732 {l}
Rbot_702_732 bot702 bot732 {r}
Lbot_702_732 bot702 bot732 {l}
C702 top702 bot702 {c}
Rtop_703_704 top703 top704 {r}
Ltop_703_704 top703 top704 {l}
Rbot_703_704 bot703 bot704 {r}
Lbot_703_704 bot703 bot704 {l}
Rtop_703_733 top703 top733 {r}
Ltop_703_733 top703 top733 {l}
Rbot_703_733 bot703 bot733 {r}
Lbot_703_733 bot703 bot733 {l}
C703 top703 bot703 {c}
Rtop_704_705 top704 top705 {r}
Ltop_704_705 top704 top705 {l}
Rbot_704_705 bot704 bot705 {r}
Lbot_704_705 bot704 bot705 {l}
Rtop_704_734 top704 top734 {r}
Ltop_704_734 top704 top734 {l}
Rbot_704_734 bot704 bot734 {r}
Lbot_704_734 bot704 bot734 {l}
C704 top704 bot704 {c}
Rtop_705_706 top705 top706 {r}
Ltop_705_706 top705 top706 {l}
Rbot_705_706 bot705 bot706 {r}
Lbot_705_706 bot705 bot706 {l}
Rtop_705_735 top705 top735 {r}
Ltop_705_735 top705 top735 {l}
Rbot_705_735 bot705 bot735 {r}
Lbot_705_735 bot705 bot735 {l}
C705 top705 bot705 {c}
Rtop_706_707 top706 top707 {r}
Ltop_706_707 top706 top707 {l}
Rbot_706_707 bot706 bot707 {r}
Lbot_706_707 bot706 bot707 {l}
Rtop_706_736 top706 top736 {r}
Ltop_706_736 top706 top736 {l}
Rbot_706_736 bot706 bot736 {r}
Lbot_706_736 bot706 bot736 {l}
C706 top706 bot706 {c}
Rtop_707_708 top707 top708 {r}
Ltop_707_708 top707 top708 {l}
Rbot_707_708 bot707 bot708 {r}
Lbot_707_708 bot707 bot708 {l}
Rtop_707_737 top707 top737 {r}
Ltop_707_737 top707 top737 {l}
Rbot_707_737 bot707 bot737 {r}
Lbot_707_737 bot707 bot737 {l}
C707 top707 bot707 {c}
Rtop_708_709 top708 top709 {r}
Ltop_708_709 top708 top709 {l}
Rbot_708_709 bot708 bot709 {r}
Lbot_708_709 bot708 bot709 {l}
Rtop_708_738 top708 top738 {r}
Ltop_708_738 top708 top738 {l}
Rbot_708_738 bot708 bot738 {r}
Lbot_708_738 bot708 bot738 {l}
C708 top708 bot708 {c}
Rtop_709_710 top709 top710 {r}
Ltop_709_710 top709 top710 {l}
Rbot_709_710 bot709 bot710 {r}
Lbot_709_710 bot709 bot710 {l}
Rtop_709_739 top709 top739 {r}
Ltop_709_739 top709 top739 {l}
Rbot_709_739 bot709 bot739 {r}
Lbot_709_739 bot709 bot739 {l}
C709 top709 bot709 {c}
Rtop_710_711 top710 top711 {r}
Ltop_710_711 top710 top711 {l}
Rbot_710_711 bot710 bot711 {r}
Lbot_710_711 bot710 bot711 {l}
Rtop_710_740 top710 top740 {r}
Ltop_710_740 top710 top740 {l}
Rbot_710_740 bot710 bot740 {r}
Lbot_710_740 bot710 bot740 {l}
C710 top710 bot710 {c}
Rtop_711_712 top711 top712 {r}
Ltop_711_712 top711 top712 {l}
Rbot_711_712 bot711 bot712 {r}
Lbot_711_712 bot711 bot712 {l}
Rtop_711_741 top711 top741 {r}
Ltop_711_741 top711 top741 {l}
Rbot_711_741 bot711 bot741 {r}
Lbot_711_741 bot711 bot741 {l}
C711 top711 bot711 {c}
Rtop_712_713 top712 top713 {r}
Ltop_712_713 top712 top713 {l}
Rbot_712_713 bot712 bot713 {r}
Lbot_712_713 bot712 bot713 {l}
Rtop_712_742 top712 top742 {r}
Ltop_712_742 top712 top742 {l}
Rbot_712_742 bot712 bot742 {r}
Lbot_712_742 bot712 bot742 {l}
C712 top712 bot712 {c}
Rtop_713_714 top713 top714 {r}
Ltop_713_714 top713 top714 {l}
Rbot_713_714 bot713 bot714 {r}
Lbot_713_714 bot713 bot714 {l}
Rtop_713_743 top713 top743 {r}
Ltop_713_743 top713 top743 {l}
Rbot_713_743 bot713 bot743 {r}
Lbot_713_743 bot713 bot743 {l}
C713 top713 bot713 {c}
Rtop_714_715 top714 top715 {r}
Ltop_714_715 top714 top715 {l}
Rbot_714_715 bot714 bot715 {r}
Lbot_714_715 bot714 bot715 {l}
Rtop_714_744 top714 top744 {r}
Ltop_714_744 top714 top744 {l}
Rbot_714_744 bot714 bot744 {r}
Lbot_714_744 bot714 bot744 {l}
C714 top714 bot714 {c}
Rtop_715_716 top715 top716 {r}
Ltop_715_716 top715 top716 {l}
Rbot_715_716 bot715 bot716 {r}
Lbot_715_716 bot715 bot716 {l}
Rtop_715_745 top715 top745 {r}
Ltop_715_745 top715 top745 {l}
Rbot_715_745 bot715 bot745 {r}
Lbot_715_745 bot715 bot745 {l}
C715 top715 bot715 {c}
Rtop_716_717 top716 top717 {r}
Ltop_716_717 top716 top717 {l}
Rbot_716_717 bot716 bot717 {r}
Lbot_716_717 bot716 bot717 {l}
Rtop_716_746 top716 top746 {r}
Ltop_716_746 top716 top746 {l}
Rbot_716_746 bot716 bot746 {r}
Lbot_716_746 bot716 bot746 {l}
C716 top716 bot716 {c}
Rtop_717_718 top717 top718 {r}
Ltop_717_718 top717 top718 {l}
Rbot_717_718 bot717 bot718 {r}
Lbot_717_718 bot717 bot718 {l}
Rtop_717_747 top717 top747 {r}
Ltop_717_747 top717 top747 {l}
Rbot_717_747 bot717 bot747 {r}
Lbot_717_747 bot717 bot747 {l}
C717 top717 bot717 {c}
Rtop_718_719 top718 top719 {r}
Ltop_718_719 top718 top719 {l}
Rbot_718_719 bot718 bot719 {r}
Lbot_718_719 bot718 bot719 {l}
Rtop_718_748 top718 top748 {r}
Ltop_718_748 top718 top748 {l}
Rbot_718_748 bot718 bot748 {r}
Lbot_718_748 bot718 bot748 {l}
C718 top718 bot718 {c}
Rtop_719_720 top719 top720 {r}
Ltop_719_720 top719 top720 {l}
Rbot_719_720 bot719 bot720 {r}
Lbot_719_720 bot719 bot720 {l}
Rtop_719_749 top719 top749 {r}
Ltop_719_749 top719 top749 {l}
Rbot_719_749 bot719 bot749 {r}
Lbot_719_749 bot719 bot749 {l}
C719 top719 bot719 {c}
Rtop_720_750 top720 top750 {r}
Ltop_720_750 top720 top750 {l}
Rbot_720_750 bot720 bot750 {r}
Lbot_720_750 bot720 bot750 {l}
C720 top720 bot720 {c}
Rtop_721_722 top721 top722 {r}
Ltop_721_722 top721 top722 {l}
Rbot_721_722 bot721 bot722 {r}
Lbot_721_722 bot721 bot722 {l}
Rtop_721_751 top721 top751 {r}
Ltop_721_751 top721 top751 {l}
Rbot_721_751 bot721 bot751 {r}
Lbot_721_751 bot721 bot751 {l}
C721 top721 bot721 {c}
Rtop_722_723 top722 top723 {r}
Ltop_722_723 top722 top723 {l}
Rbot_722_723 bot722 bot723 {r}
Lbot_722_723 bot722 bot723 {l}
Rtop_722_752 top722 top752 {r}
Ltop_722_752 top722 top752 {l}
Rbot_722_752 bot722 bot752 {r}
Lbot_722_752 bot722 bot752 {l}
C722 top722 bot722 {c}
Rtop_723_724 top723 top724 {r}
Ltop_723_724 top723 top724 {l}
Rbot_723_724 bot723 bot724 {r}
Lbot_723_724 bot723 bot724 {l}
Rtop_723_753 top723 top753 {r}
Ltop_723_753 top723 top753 {l}
Rbot_723_753 bot723 bot753 {r}
Lbot_723_753 bot723 bot753 {l}
C723 top723 bot723 {c}
Rtop_724_725 top724 top725 {r}
Ltop_724_725 top724 top725 {l}
Rbot_724_725 bot724 bot725 {r}
Lbot_724_725 bot724 bot725 {l}
Rtop_724_754 top724 top754 {r}
Ltop_724_754 top724 top754 {l}
Rbot_724_754 bot724 bot754 {r}
Lbot_724_754 bot724 bot754 {l}
C724 top724 bot724 {c}
Rtop_725_726 top725 top726 {r}
Ltop_725_726 top725 top726 {l}
Rbot_725_726 bot725 bot726 {r}
Lbot_725_726 bot725 bot726 {l}
Rtop_725_755 top725 top755 {r}
Ltop_725_755 top725 top755 {l}
Rbot_725_755 bot725 bot755 {r}
Lbot_725_755 bot725 bot755 {l}
C725 top725 bot725 {c}
Rtop_726_727 top726 top727 {r}
Ltop_726_727 top726 top727 {l}
Rbot_726_727 bot726 bot727 {r}
Lbot_726_727 bot726 bot727 {l}
Rtop_726_756 top726 top756 {r}
Ltop_726_756 top726 top756 {l}
Rbot_726_756 bot726 bot756 {r}
Lbot_726_756 bot726 bot756 {l}
C726 top726 bot726 {c}
Rtop_727_728 top727 top728 {r}
Ltop_727_728 top727 top728 {l}
Rbot_727_728 bot727 bot728 {r}
Lbot_727_728 bot727 bot728 {l}
Rtop_727_757 top727 top757 {r}
Ltop_727_757 top727 top757 {l}
Rbot_727_757 bot727 bot757 {r}
Lbot_727_757 bot727 bot757 {l}
C727 top727 bot727 {c}
Rtop_728_729 top728 top729 {r}
Ltop_728_729 top728 top729 {l}
Rbot_728_729 bot728 bot729 {r}
Lbot_728_729 bot728 bot729 {l}
Rtop_728_758 top728 top758 {r}
Ltop_728_758 top728 top758 {l}
Rbot_728_758 bot728 bot758 {r}
Lbot_728_758 bot728 bot758 {l}
C728 top728 bot728 {c}
Rtop_729_730 top729 top730 {r}
Ltop_729_730 top729 top730 {l}
Rbot_729_730 bot729 bot730 {r}
Lbot_729_730 bot729 bot730 {l}
Rtop_729_759 top729 top759 {r}
Ltop_729_759 top729 top759 {l}
Rbot_729_759 bot729 bot759 {r}
Lbot_729_759 bot729 bot759 {l}
C729 top729 bot729 {c}
Rtop_730_731 top730 top731 {r}
Ltop_730_731 top730 top731 {l}
Rbot_730_731 bot730 bot731 {r}
Lbot_730_731 bot730 bot731 {l}
Rtop_730_760 top730 top760 {r}
Ltop_730_760 top730 top760 {l}
Rbot_730_760 bot730 bot760 {r}
Lbot_730_760 bot730 bot760 {l}
C730 top730 bot730 {c}
Rtop_731_732 top731 top732 {r}
Ltop_731_732 top731 top732 {l}
Rbot_731_732 bot731 bot732 {r}
Lbot_731_732 bot731 bot732 {l}
Rtop_731_761 top731 top761 {r}
Ltop_731_761 top731 top761 {l}
Rbot_731_761 bot731 bot761 {r}
Lbot_731_761 bot731 bot761 {l}
C731 top731 bot731 {c}
Rtop_732_733 top732 top733 {r}
Ltop_732_733 top732 top733 {l}
Rbot_732_733 bot732 bot733 {r}
Lbot_732_733 bot732 bot733 {l}
Rtop_732_762 top732 top762 {r}
Ltop_732_762 top732 top762 {l}
Rbot_732_762 bot732 bot762 {r}
Lbot_732_762 bot732 bot762 {l}
C732 top732 bot732 {c}
Rtop_733_734 top733 top734 {r}
Ltop_733_734 top733 top734 {l}
Rbot_733_734 bot733 bot734 {r}
Lbot_733_734 bot733 bot734 {l}
Rtop_733_763 top733 top763 {r}
Ltop_733_763 top733 top763 {l}
Rbot_733_763 bot733 bot763 {r}
Lbot_733_763 bot733 bot763 {l}
C733 top733 bot733 {c}
Rtop_734_735 top734 top735 {r}
Ltop_734_735 top734 top735 {l}
Rbot_734_735 bot734 bot735 {r}
Lbot_734_735 bot734 bot735 {l}
Rtop_734_764 top734 top764 {r}
Ltop_734_764 top734 top764 {l}
Rbot_734_764 bot734 bot764 {r}
Lbot_734_764 bot734 bot764 {l}
C734 top734 bot734 {c}
Rtop_735_736 top735 top736 {r}
Ltop_735_736 top735 top736 {l}
Rbot_735_736 bot735 bot736 {r}
Lbot_735_736 bot735 bot736 {l}
Rtop_735_765 top735 top765 {r}
Ltop_735_765 top735 top765 {l}
Rbot_735_765 bot735 bot765 {r}
Lbot_735_765 bot735 bot765 {l}
C735 top735 bot735 {c}
Rtop_736_737 top736 top737 {r}
Ltop_736_737 top736 top737 {l}
Rbot_736_737 bot736 bot737 {r}
Lbot_736_737 bot736 bot737 {l}
Rtop_736_766 top736 top766 {r}
Ltop_736_766 top736 top766 {l}
Rbot_736_766 bot736 bot766 {r}
Lbot_736_766 bot736 bot766 {l}
C736 top736 bot736 {c}
Rtop_737_738 top737 top738 {r}
Ltop_737_738 top737 top738 {l}
Rbot_737_738 bot737 bot738 {r}
Lbot_737_738 bot737 bot738 {l}
Rtop_737_767 top737 top767 {r}
Ltop_737_767 top737 top767 {l}
Rbot_737_767 bot737 bot767 {r}
Lbot_737_767 bot737 bot767 {l}
C737 top737 bot737 {c}
Rtop_738_739 top738 top739 {r}
Ltop_738_739 top738 top739 {l}
Rbot_738_739 bot738 bot739 {r}
Lbot_738_739 bot738 bot739 {l}
Rtop_738_768 top738 top768 {r}
Ltop_738_768 top738 top768 {l}
Rbot_738_768 bot738 bot768 {r}
Lbot_738_768 bot738 bot768 {l}
C738 top738 bot738 {c}
Rtop_739_740 top739 top740 {r}
Ltop_739_740 top739 top740 {l}
Rbot_739_740 bot739 bot740 {r}
Lbot_739_740 bot739 bot740 {l}
Rtop_739_769 top739 top769 {r}
Ltop_739_769 top739 top769 {l}
Rbot_739_769 bot739 bot769 {r}
Lbot_739_769 bot739 bot769 {l}
C739 top739 bot739 {c}
Rtop_740_741 top740 top741 {r}
Ltop_740_741 top740 top741 {l}
Rbot_740_741 bot740 bot741 {r}
Lbot_740_741 bot740 bot741 {l}
Rtop_740_770 top740 top770 {r}
Ltop_740_770 top740 top770 {l}
Rbot_740_770 bot740 bot770 {r}
Lbot_740_770 bot740 bot770 {l}
C740 top740 bot740 {c}
Rtop_741_742 top741 top742 {r}
Ltop_741_742 top741 top742 {l}
Rbot_741_742 bot741 bot742 {r}
Lbot_741_742 bot741 bot742 {l}
Rtop_741_771 top741 top771 {r}
Ltop_741_771 top741 top771 {l}
Rbot_741_771 bot741 bot771 {r}
Lbot_741_771 bot741 bot771 {l}
C741 top741 bot741 {c}
Rtop_742_743 top742 top743 {r}
Ltop_742_743 top742 top743 {l}
Rbot_742_743 bot742 bot743 {r}
Lbot_742_743 bot742 bot743 {l}
Rtop_742_772 top742 top772 {r}
Ltop_742_772 top742 top772 {l}
Rbot_742_772 bot742 bot772 {r}
Lbot_742_772 bot742 bot772 {l}
C742 top742 bot742 {c}
Rtop_743_744 top743 top744 {r}
Ltop_743_744 top743 top744 {l}
Rbot_743_744 bot743 bot744 {r}
Lbot_743_744 bot743 bot744 {l}
Rtop_743_773 top743 top773 {r}
Ltop_743_773 top743 top773 {l}
Rbot_743_773 bot743 bot773 {r}
Lbot_743_773 bot743 bot773 {l}
C743 top743 bot743 {c}
Rtop_744_745 top744 top745 {r}
Ltop_744_745 top744 top745 {l}
Rbot_744_745 bot744 bot745 {r}
Lbot_744_745 bot744 bot745 {l}
Rtop_744_774 top744 top774 {r}
Ltop_744_774 top744 top774 {l}
Rbot_744_774 bot744 bot774 {r}
Lbot_744_774 bot744 bot774 {l}
C744 top744 bot744 {c}
Rtop_745_746 top745 top746 {r}
Ltop_745_746 top745 top746 {l}
Rbot_745_746 bot745 bot746 {r}
Lbot_745_746 bot745 bot746 {l}
Rtop_745_775 top745 top775 {r}
Ltop_745_775 top745 top775 {l}
Rbot_745_775 bot745 bot775 {r}
Lbot_745_775 bot745 bot775 {l}
C745 top745 bot745 {c}
Rtop_746_747 top746 top747 {r}
Ltop_746_747 top746 top747 {l}
Rbot_746_747 bot746 bot747 {r}
Lbot_746_747 bot746 bot747 {l}
Rtop_746_776 top746 top776 {r}
Ltop_746_776 top746 top776 {l}
Rbot_746_776 bot746 bot776 {r}
Lbot_746_776 bot746 bot776 {l}
C746 top746 bot746 {c}
Rtop_747_748 top747 top748 {r}
Ltop_747_748 top747 top748 {l}
Rbot_747_748 bot747 bot748 {r}
Lbot_747_748 bot747 bot748 {l}
Rtop_747_777 top747 top777 {r}
Ltop_747_777 top747 top777 {l}
Rbot_747_777 bot747 bot777 {r}
Lbot_747_777 bot747 bot777 {l}
C747 top747 bot747 {c}
Rtop_748_749 top748 top749 {r}
Ltop_748_749 top748 top749 {l}
Rbot_748_749 bot748 bot749 {r}
Lbot_748_749 bot748 bot749 {l}
Rtop_748_778 top748 top778 {r}
Ltop_748_778 top748 top778 {l}
Rbot_748_778 bot748 bot778 {r}
Lbot_748_778 bot748 bot778 {l}
C748 top748 bot748 {c}
Rtop_749_750 top749 top750 {r}
Ltop_749_750 top749 top750 {l}
Rbot_749_750 bot749 bot750 {r}
Lbot_749_750 bot749 bot750 {l}
Rtop_749_779 top749 top779 {r}
Ltop_749_779 top749 top779 {l}
Rbot_749_779 bot749 bot779 {r}
Lbot_749_779 bot749 bot779 {l}
C749 top749 bot749 {c}
Rtop_750_780 top750 top780 {r}
Ltop_750_780 top750 top780 {l}
Rbot_750_780 bot750 bot780 {r}
Lbot_750_780 bot750 bot780 {l}
C750 top750 bot750 {c}
Rtop_751_752 top751 top752 {r}
Ltop_751_752 top751 top752 {l}
Rbot_751_752 bot751 bot752 {r}
Lbot_751_752 bot751 bot752 {l}
Rtop_751_781 top751 top781 {r}
Ltop_751_781 top751 top781 {l}
Rbot_751_781 bot751 bot781 {r}
Lbot_751_781 bot751 bot781 {l}
C751 top751 bot751 {c}
Rtop_752_753 top752 top753 {r}
Ltop_752_753 top752 top753 {l}
Rbot_752_753 bot752 bot753 {r}
Lbot_752_753 bot752 bot753 {l}
Rtop_752_782 top752 top782 {r}
Ltop_752_782 top752 top782 {l}
Rbot_752_782 bot752 bot782 {r}
Lbot_752_782 bot752 bot782 {l}
C752 top752 bot752 {c}
Rtop_753_754 top753 top754 {r}
Ltop_753_754 top753 top754 {l}
Rbot_753_754 bot753 bot754 {r}
Lbot_753_754 bot753 bot754 {l}
Rtop_753_783 top753 top783 {r}
Ltop_753_783 top753 top783 {l}
Rbot_753_783 bot753 bot783 {r}
Lbot_753_783 bot753 bot783 {l}
C753 top753 bot753 {c}
Rtop_754_755 top754 top755 {r}
Ltop_754_755 top754 top755 {l}
Rbot_754_755 bot754 bot755 {r}
Lbot_754_755 bot754 bot755 {l}
Rtop_754_784 top754 top784 {r}
Ltop_754_784 top754 top784 {l}
Rbot_754_784 bot754 bot784 {r}
Lbot_754_784 bot754 bot784 {l}
C754 top754 bot754 {c}
Rtop_755_756 top755 top756 {r}
Ltop_755_756 top755 top756 {l}
Rbot_755_756 bot755 bot756 {r}
Lbot_755_756 bot755 bot756 {l}
Rtop_755_785 top755 top785 {r}
Ltop_755_785 top755 top785 {l}
Rbot_755_785 bot755 bot785 {r}
Lbot_755_785 bot755 bot785 {l}
C755 top755 bot755 {c}
Rtop_756_757 top756 top757 {r}
Ltop_756_757 top756 top757 {l}
Rbot_756_757 bot756 bot757 {r}
Lbot_756_757 bot756 bot757 {l}
Rtop_756_786 top756 top786 {r}
Ltop_756_786 top756 top786 {l}
Rbot_756_786 bot756 bot786 {r}
Lbot_756_786 bot756 bot786 {l}
C756 top756 bot756 {c}
Rtop_757_758 top757 top758 {r}
Ltop_757_758 top757 top758 {l}
Rbot_757_758 bot757 bot758 {r}
Lbot_757_758 bot757 bot758 {l}
Rtop_757_787 top757 top787 {r}
Ltop_757_787 top757 top787 {l}
Rbot_757_787 bot757 bot787 {r}
Lbot_757_787 bot757 bot787 {l}
C757 top757 bot757 {c}
Rtop_758_759 top758 top759 {r}
Ltop_758_759 top758 top759 {l}
Rbot_758_759 bot758 bot759 {r}
Lbot_758_759 bot758 bot759 {l}
Rtop_758_788 top758 top788 {r}
Ltop_758_788 top758 top788 {l}
Rbot_758_788 bot758 bot788 {r}
Lbot_758_788 bot758 bot788 {l}
C758 top758 bot758 {c}
Rtop_759_760 top759 top760 {r}
Ltop_759_760 top759 top760 {l}
Rbot_759_760 bot759 bot760 {r}
Lbot_759_760 bot759 bot760 {l}
Rtop_759_789 top759 top789 {r}
Ltop_759_789 top759 top789 {l}
Rbot_759_789 bot759 bot789 {r}
Lbot_759_789 bot759 bot789 {l}
C759 top759 bot759 {c}
Rtop_760_761 top760 top761 {r}
Ltop_760_761 top760 top761 {l}
Rbot_760_761 bot760 bot761 {r}
Lbot_760_761 bot760 bot761 {l}
Rtop_760_790 top760 top790 {r}
Ltop_760_790 top760 top790 {l}
Rbot_760_790 bot760 bot790 {r}
Lbot_760_790 bot760 bot790 {l}
C760 top760 bot760 {c}
Rtop_761_762 top761 top762 {r}
Ltop_761_762 top761 top762 {l}
Rbot_761_762 bot761 bot762 {r}
Lbot_761_762 bot761 bot762 {l}
Rtop_761_791 top761 top791 {r}
Ltop_761_791 top761 top791 {l}
Rbot_761_791 bot761 bot791 {r}
Lbot_761_791 bot761 bot791 {l}
C761 top761 bot761 {c}
Rtop_762_763 top762 top763 {r}
Ltop_762_763 top762 top763 {l}
Rbot_762_763 bot762 bot763 {r}
Lbot_762_763 bot762 bot763 {l}
Rtop_762_792 top762 top792 {r}
Ltop_762_792 top762 top792 {l}
Rbot_762_792 bot762 bot792 {r}
Lbot_762_792 bot762 bot792 {l}
C762 top762 bot762 {c}
Rtop_763_764 top763 top764 {r}
Ltop_763_764 top763 top764 {l}
Rbot_763_764 bot763 bot764 {r}
Lbot_763_764 bot763 bot764 {l}
Rtop_763_793 top763 top793 {r}
Ltop_763_793 top763 top793 {l}
Rbot_763_793 bot763 bot793 {r}
Lbot_763_793 bot763 bot793 {l}
C763 top763 bot763 {c}
Rtop_764_765 top764 top765 {r}
Ltop_764_765 top764 top765 {l}
Rbot_764_765 bot764 bot765 {r}
Lbot_764_765 bot764 bot765 {l}
Rtop_764_794 top764 top794 {r}
Ltop_764_794 top764 top794 {l}
Rbot_764_794 bot764 bot794 {r}
Lbot_764_794 bot764 bot794 {l}
C764 top764 bot764 {c}
Rtop_765_766 top765 top766 {r}
Ltop_765_766 top765 top766 {l}
Rbot_765_766 bot765 bot766 {r}
Lbot_765_766 bot765 bot766 {l}
Rtop_765_795 top765 top795 {r}
Ltop_765_795 top765 top795 {l}
Rbot_765_795 bot765 bot795 {r}
Lbot_765_795 bot765 bot795 {l}
C765 top765 bot765 {c}
Rtop_766_767 top766 top767 {r}
Ltop_766_767 top766 top767 {l}
Rbot_766_767 bot766 bot767 {r}
Lbot_766_767 bot766 bot767 {l}
Rtop_766_796 top766 top796 {r}
Ltop_766_796 top766 top796 {l}
Rbot_766_796 bot766 bot796 {r}
Lbot_766_796 bot766 bot796 {l}
C766 top766 bot766 {c}
Rtop_767_768 top767 top768 {r}
Ltop_767_768 top767 top768 {l}
Rbot_767_768 bot767 bot768 {r}
Lbot_767_768 bot767 bot768 {l}
Rtop_767_797 top767 top797 {r}
Ltop_767_797 top767 top797 {l}
Rbot_767_797 bot767 bot797 {r}
Lbot_767_797 bot767 bot797 {l}
C767 top767 bot767 {c}
Rtop_768_769 top768 top769 {r}
Ltop_768_769 top768 top769 {l}
Rbot_768_769 bot768 bot769 {r}
Lbot_768_769 bot768 bot769 {l}
Rtop_768_798 top768 top798 {r}
Ltop_768_798 top768 top798 {l}
Rbot_768_798 bot768 bot798 {r}
Lbot_768_798 bot768 bot798 {l}
C768 top768 bot768 {c}
Rtop_769_770 top769 top770 {r}
Ltop_769_770 top769 top770 {l}
Rbot_769_770 bot769 bot770 {r}
Lbot_769_770 bot769 bot770 {l}
Rtop_769_799 top769 top799 {r}
Ltop_769_799 top769 top799 {l}
Rbot_769_799 bot769 bot799 {r}
Lbot_769_799 bot769 bot799 {l}
C769 top769 bot769 {c}
Rtop_770_771 top770 top771 {r}
Ltop_770_771 top770 top771 {l}
Rbot_770_771 bot770 bot771 {r}
Lbot_770_771 bot770 bot771 {l}
Rtop_770_800 top770 top800 {r}
Ltop_770_800 top770 top800 {l}
Rbot_770_800 bot770 bot800 {r}
Lbot_770_800 bot770 bot800 {l}
C770 top770 bot770 {c}
Rtop_771_772 top771 top772 {r}
Ltop_771_772 top771 top772 {l}
Rbot_771_772 bot771 bot772 {r}
Lbot_771_772 bot771 bot772 {l}
Rtop_771_801 top771 top801 {r}
Ltop_771_801 top771 top801 {l}
Rbot_771_801 bot771 bot801 {r}
Lbot_771_801 bot771 bot801 {l}
C771 top771 bot771 {c}
Rtop_772_773 top772 top773 {r}
Ltop_772_773 top772 top773 {l}
Rbot_772_773 bot772 bot773 {r}
Lbot_772_773 bot772 bot773 {l}
Rtop_772_802 top772 top802 {r}
Ltop_772_802 top772 top802 {l}
Rbot_772_802 bot772 bot802 {r}
Lbot_772_802 bot772 bot802 {l}
C772 top772 bot772 {c}
Rtop_773_774 top773 top774 {r}
Ltop_773_774 top773 top774 {l}
Rbot_773_774 bot773 bot774 {r}
Lbot_773_774 bot773 bot774 {l}
Rtop_773_803 top773 top803 {r}
Ltop_773_803 top773 top803 {l}
Rbot_773_803 bot773 bot803 {r}
Lbot_773_803 bot773 bot803 {l}
C773 top773 bot773 {c}
Rtop_774_775 top774 top775 {r}
Ltop_774_775 top774 top775 {l}
Rbot_774_775 bot774 bot775 {r}
Lbot_774_775 bot774 bot775 {l}
Rtop_774_804 top774 top804 {r}
Ltop_774_804 top774 top804 {l}
Rbot_774_804 bot774 bot804 {r}
Lbot_774_804 bot774 bot804 {l}
C774 top774 bot774 {c}
Rtop_775_776 top775 top776 {r}
Ltop_775_776 top775 top776 {l}
Rbot_775_776 bot775 bot776 {r}
Lbot_775_776 bot775 bot776 {l}
Rtop_775_805 top775 top805 {r}
Ltop_775_805 top775 top805 {l}
Rbot_775_805 bot775 bot805 {r}
Lbot_775_805 bot775 bot805 {l}
C775 top775 bot775 {c}
Rtop_776_777 top776 top777 {r}
Ltop_776_777 top776 top777 {l}
Rbot_776_777 bot776 bot777 {r}
Lbot_776_777 bot776 bot777 {l}
Rtop_776_806 top776 top806 {r}
Ltop_776_806 top776 top806 {l}
Rbot_776_806 bot776 bot806 {r}
Lbot_776_806 bot776 bot806 {l}
C776 top776 bot776 {c}
Rtop_777_778 top777 top778 {r}
Ltop_777_778 top777 top778 {l}
Rbot_777_778 bot777 bot778 {r}
Lbot_777_778 bot777 bot778 {l}
Rtop_777_807 top777 top807 {r}
Ltop_777_807 top777 top807 {l}
Rbot_777_807 bot777 bot807 {r}
Lbot_777_807 bot777 bot807 {l}
C777 top777 bot777 {c}
Rtop_778_779 top778 top779 {r}
Ltop_778_779 top778 top779 {l}
Rbot_778_779 bot778 bot779 {r}
Lbot_778_779 bot778 bot779 {l}
Rtop_778_808 top778 top808 {r}
Ltop_778_808 top778 top808 {l}
Rbot_778_808 bot778 bot808 {r}
Lbot_778_808 bot778 bot808 {l}
C778 top778 bot778 {c}
Rtop_779_780 top779 top780 {r}
Ltop_779_780 top779 top780 {l}
Rbot_779_780 bot779 bot780 {r}
Lbot_779_780 bot779 bot780 {l}
Rtop_779_809 top779 top809 {r}
Ltop_779_809 top779 top809 {l}
Rbot_779_809 bot779 bot809 {r}
Lbot_779_809 bot779 bot809 {l}
C779 top779 bot779 {c}
Rtop_780_810 top780 top810 {r}
Ltop_780_810 top780 top810 {l}
Rbot_780_810 bot780 bot810 {r}
Lbot_780_810 bot780 bot810 {l}
C780 top780 bot780 {c}
Rtop_781_782 top781 top782 {r}
Ltop_781_782 top781 top782 {l}
Rbot_781_782 bot781 bot782 {r}
Lbot_781_782 bot781 bot782 {l}
Rtop_781_811 top781 top811 {r}
Ltop_781_811 top781 top811 {l}
Rbot_781_811 bot781 bot811 {r}
Lbot_781_811 bot781 bot811 {l}
C781 top781 bot781 {c}
Rtop_782_783 top782 top783 {r}
Ltop_782_783 top782 top783 {l}
Rbot_782_783 bot782 bot783 {r}
Lbot_782_783 bot782 bot783 {l}
Rtop_782_812 top782 top812 {r}
Ltop_782_812 top782 top812 {l}
Rbot_782_812 bot782 bot812 {r}
Lbot_782_812 bot782 bot812 {l}
C782 top782 bot782 {c}
Rtop_783_784 top783 top784 {r}
Ltop_783_784 top783 top784 {l}
Rbot_783_784 bot783 bot784 {r}
Lbot_783_784 bot783 bot784 {l}
Rtop_783_813 top783 top813 {r}
Ltop_783_813 top783 top813 {l}
Rbot_783_813 bot783 bot813 {r}
Lbot_783_813 bot783 bot813 {l}
C783 top783 bot783 {c}
Rtop_784_785 top784 top785 {r}
Ltop_784_785 top784 top785 {l}
Rbot_784_785 bot784 bot785 {r}
Lbot_784_785 bot784 bot785 {l}
Rtop_784_814 top784 top814 {r}
Ltop_784_814 top784 top814 {l}
Rbot_784_814 bot784 bot814 {r}
Lbot_784_814 bot784 bot814 {l}
C784 top784 bot784 {c}
Rtop_785_786 top785 top786 {r}
Ltop_785_786 top785 top786 {l}
Rbot_785_786 bot785 bot786 {r}
Lbot_785_786 bot785 bot786 {l}
Rtop_785_815 top785 top815 {r}
Ltop_785_815 top785 top815 {l}
Rbot_785_815 bot785 bot815 {r}
Lbot_785_815 bot785 bot815 {l}
C785 top785 bot785 {c}
Rtop_786_787 top786 top787 {r}
Ltop_786_787 top786 top787 {l}
Rbot_786_787 bot786 bot787 {r}
Lbot_786_787 bot786 bot787 {l}
Rtop_786_816 top786 top816 {r}
Ltop_786_816 top786 top816 {l}
Rbot_786_816 bot786 bot816 {r}
Lbot_786_816 bot786 bot816 {l}
C786 top786 bot786 {c}
Rtop_787_788 top787 top788 {r}
Ltop_787_788 top787 top788 {l}
Rbot_787_788 bot787 bot788 {r}
Lbot_787_788 bot787 bot788 {l}
Rtop_787_817 top787 top817 {r}
Ltop_787_817 top787 top817 {l}
Rbot_787_817 bot787 bot817 {r}
Lbot_787_817 bot787 bot817 {l}
C787 top787 bot787 {c}
Rtop_788_789 top788 top789 {r}
Ltop_788_789 top788 top789 {l}
Rbot_788_789 bot788 bot789 {r}
Lbot_788_789 bot788 bot789 {l}
Rtop_788_818 top788 top818 {r}
Ltop_788_818 top788 top818 {l}
Rbot_788_818 bot788 bot818 {r}
Lbot_788_818 bot788 bot818 {l}
C788 top788 bot788 {c}
Rtop_789_790 top789 top790 {r}
Ltop_789_790 top789 top790 {l}
Rbot_789_790 bot789 bot790 {r}
Lbot_789_790 bot789 bot790 {l}
Rtop_789_819 top789 top819 {r}
Ltop_789_819 top789 top819 {l}
Rbot_789_819 bot789 bot819 {r}
Lbot_789_819 bot789 bot819 {l}
C789 top789 bot789 {c}
Rtop_790_791 top790 top791 {r}
Ltop_790_791 top790 top791 {l}
Rbot_790_791 bot790 bot791 {r}
Lbot_790_791 bot790 bot791 {l}
Rtop_790_820 top790 top820 {r}
Ltop_790_820 top790 top820 {l}
Rbot_790_820 bot790 bot820 {r}
Lbot_790_820 bot790 bot820 {l}
C790 top790 bot790 {c}
Rtop_791_792 top791 top792 {r}
Ltop_791_792 top791 top792 {l}
Rbot_791_792 bot791 bot792 {r}
Lbot_791_792 bot791 bot792 {l}
Rtop_791_821 top791 top821 {r}
Ltop_791_821 top791 top821 {l}
Rbot_791_821 bot791 bot821 {r}
Lbot_791_821 bot791 bot821 {l}
C791 top791 bot791 {c}
Rtop_792_793 top792 top793 {r}
Ltop_792_793 top792 top793 {l}
Rbot_792_793 bot792 bot793 {r}
Lbot_792_793 bot792 bot793 {l}
Rtop_792_822 top792 top822 {r}
Ltop_792_822 top792 top822 {l}
Rbot_792_822 bot792 bot822 {r}
Lbot_792_822 bot792 bot822 {l}
C792 top792 bot792 {c}
Rtop_793_794 top793 top794 {r}
Ltop_793_794 top793 top794 {l}
Rbot_793_794 bot793 bot794 {r}
Lbot_793_794 bot793 bot794 {l}
Rtop_793_823 top793 top823 {r}
Ltop_793_823 top793 top823 {l}
Rbot_793_823 bot793 bot823 {r}
Lbot_793_823 bot793 bot823 {l}
C793 top793 bot793 {c}
Rtop_794_795 top794 top795 {r}
Ltop_794_795 top794 top795 {l}
Rbot_794_795 bot794 bot795 {r}
Lbot_794_795 bot794 bot795 {l}
Rtop_794_824 top794 top824 {r}
Ltop_794_824 top794 top824 {l}
Rbot_794_824 bot794 bot824 {r}
Lbot_794_824 bot794 bot824 {l}
C794 top794 bot794 {c}
Rtop_795_796 top795 top796 {r}
Ltop_795_796 top795 top796 {l}
Rbot_795_796 bot795 bot796 {r}
Lbot_795_796 bot795 bot796 {l}
Rtop_795_825 top795 top825 {r}
Ltop_795_825 top795 top825 {l}
Rbot_795_825 bot795 bot825 {r}
Lbot_795_825 bot795 bot825 {l}
C795 top795 bot795 {c}
Rtop_796_797 top796 top797 {r}
Ltop_796_797 top796 top797 {l}
Rbot_796_797 bot796 bot797 {r}
Lbot_796_797 bot796 bot797 {l}
Rtop_796_826 top796 top826 {r}
Ltop_796_826 top796 top826 {l}
Rbot_796_826 bot796 bot826 {r}
Lbot_796_826 bot796 bot826 {l}
C796 top796 bot796 {c}
Rtop_797_798 top797 top798 {r}
Ltop_797_798 top797 top798 {l}
Rbot_797_798 bot797 bot798 {r}
Lbot_797_798 bot797 bot798 {l}
Rtop_797_827 top797 top827 {r}
Ltop_797_827 top797 top827 {l}
Rbot_797_827 bot797 bot827 {r}
Lbot_797_827 bot797 bot827 {l}
C797 top797 bot797 {c}
Rtop_798_799 top798 top799 {r}
Ltop_798_799 top798 top799 {l}
Rbot_798_799 bot798 bot799 {r}
Lbot_798_799 bot798 bot799 {l}
Rtop_798_828 top798 top828 {r}
Ltop_798_828 top798 top828 {l}
Rbot_798_828 bot798 bot828 {r}
Lbot_798_828 bot798 bot828 {l}
C798 top798 bot798 {c}
Rtop_799_800 top799 top800 {r}
Ltop_799_800 top799 top800 {l}
Rbot_799_800 bot799 bot800 {r}
Lbot_799_800 bot799 bot800 {l}
Rtop_799_829 top799 top829 {r}
Ltop_799_829 top799 top829 {l}
Rbot_799_829 bot799 bot829 {r}
Lbot_799_829 bot799 bot829 {l}
C799 top799 bot799 {c}
Rtop_800_801 top800 top801 {r}
Ltop_800_801 top800 top801 {l}
Rbot_800_801 bot800 bot801 {r}
Lbot_800_801 bot800 bot801 {l}
Rtop_800_830 top800 top830 {r}
Ltop_800_830 top800 top830 {l}
Rbot_800_830 bot800 bot830 {r}
Lbot_800_830 bot800 bot830 {l}
C800 top800 bot800 {c}
Rtop_801_802 top801 top802 {r}
Ltop_801_802 top801 top802 {l}
Rbot_801_802 bot801 bot802 {r}
Lbot_801_802 bot801 bot802 {l}
Rtop_801_831 top801 top831 {r}
Ltop_801_831 top801 top831 {l}
Rbot_801_831 bot801 bot831 {r}
Lbot_801_831 bot801 bot831 {l}
C801 top801 bot801 {c}
Rtop_802_803 top802 top803 {r}
Ltop_802_803 top802 top803 {l}
Rbot_802_803 bot802 bot803 {r}
Lbot_802_803 bot802 bot803 {l}
Rtop_802_832 top802 top832 {r}
Ltop_802_832 top802 top832 {l}
Rbot_802_832 bot802 bot832 {r}
Lbot_802_832 bot802 bot832 {l}
C802 top802 bot802 {c}
Rtop_803_804 top803 top804 {r}
Ltop_803_804 top803 top804 {l}
Rbot_803_804 bot803 bot804 {r}
Lbot_803_804 bot803 bot804 {l}
Rtop_803_833 top803 top833 {r}
Ltop_803_833 top803 top833 {l}
Rbot_803_833 bot803 bot833 {r}
Lbot_803_833 bot803 bot833 {l}
C803 top803 bot803 {c}
Rtop_804_805 top804 top805 {r}
Ltop_804_805 top804 top805 {l}
Rbot_804_805 bot804 bot805 {r}
Lbot_804_805 bot804 bot805 {l}
Rtop_804_834 top804 top834 {r}
Ltop_804_834 top804 top834 {l}
Rbot_804_834 bot804 bot834 {r}
Lbot_804_834 bot804 bot834 {l}
C804 top804 bot804 {c}
Rtop_805_806 top805 top806 {r}
Ltop_805_806 top805 top806 {l}
Rbot_805_806 bot805 bot806 {r}
Lbot_805_806 bot805 bot806 {l}
Rtop_805_835 top805 top835 {r}
Ltop_805_835 top805 top835 {l}
Rbot_805_835 bot805 bot835 {r}
Lbot_805_835 bot805 bot835 {l}
C805 top805 bot805 {c}
Rtop_806_807 top806 top807 {r}
Ltop_806_807 top806 top807 {l}
Rbot_806_807 bot806 bot807 {r}
Lbot_806_807 bot806 bot807 {l}
Rtop_806_836 top806 top836 {r}
Ltop_806_836 top806 top836 {l}
Rbot_806_836 bot806 bot836 {r}
Lbot_806_836 bot806 bot836 {l}
C806 top806 bot806 {c}
Rtop_807_808 top807 top808 {r}
Ltop_807_808 top807 top808 {l}
Rbot_807_808 bot807 bot808 {r}
Lbot_807_808 bot807 bot808 {l}
Rtop_807_837 top807 top837 {r}
Ltop_807_837 top807 top837 {l}
Rbot_807_837 bot807 bot837 {r}
Lbot_807_837 bot807 bot837 {l}
C807 top807 bot807 {c}
Rtop_808_809 top808 top809 {r}
Ltop_808_809 top808 top809 {l}
Rbot_808_809 bot808 bot809 {r}
Lbot_808_809 bot808 bot809 {l}
Rtop_808_838 top808 top838 {r}
Ltop_808_838 top808 top838 {l}
Rbot_808_838 bot808 bot838 {r}
Lbot_808_838 bot808 bot838 {l}
C808 top808 bot808 {c}
Rtop_809_810 top809 top810 {r}
Ltop_809_810 top809 top810 {l}
Rbot_809_810 bot809 bot810 {r}
Lbot_809_810 bot809 bot810 {l}
Rtop_809_839 top809 top839 {r}
Ltop_809_839 top809 top839 {l}
Rbot_809_839 bot809 bot839 {r}
Lbot_809_839 bot809 bot839 {l}
C809 top809 bot809 {c}
Rtop_810_840 top810 top840 {r}
Ltop_810_840 top810 top840 {l}
Rbot_810_840 bot810 bot840 {r}
Lbot_810_840 bot810 bot840 {l}
C810 top810 bot810 {c}
Rtop_811_812 top811 top812 {r}
Ltop_811_812 top811 top812 {l}
Rbot_811_812 bot811 bot812 {r}
Lbot_811_812 bot811 bot812 {l}
Rtop_811_841 top811 top841 {r}
Ltop_811_841 top811 top841 {l}
Rbot_811_841 bot811 bot841 {r}
Lbot_811_841 bot811 bot841 {l}
C811 top811 bot811 {c}
Rtop_812_813 top812 top813 {r}
Ltop_812_813 top812 top813 {l}
Rbot_812_813 bot812 bot813 {r}
Lbot_812_813 bot812 bot813 {l}
Rtop_812_842 top812 top842 {r}
Ltop_812_842 top812 top842 {l}
Rbot_812_842 bot812 bot842 {r}
Lbot_812_842 bot812 bot842 {l}
C812 top812 bot812 {c}
Rtop_813_814 top813 top814 {r}
Ltop_813_814 top813 top814 {l}
Rbot_813_814 bot813 bot814 {r}
Lbot_813_814 bot813 bot814 {l}
Rtop_813_843 top813 top843 {r}
Ltop_813_843 top813 top843 {l}
Rbot_813_843 bot813 bot843 {r}
Lbot_813_843 bot813 bot843 {l}
C813 top813 bot813 {c}
Rtop_814_815 top814 top815 {r}
Ltop_814_815 top814 top815 {l}
Rbot_814_815 bot814 bot815 {r}
Lbot_814_815 bot814 bot815 {l}
Rtop_814_844 top814 top844 {r}
Ltop_814_844 top814 top844 {l}
Rbot_814_844 bot814 bot844 {r}
Lbot_814_844 bot814 bot844 {l}
C814 top814 bot814 {c}
Rtop_815_816 top815 top816 {r}
Ltop_815_816 top815 top816 {l}
Rbot_815_816 bot815 bot816 {r}
Lbot_815_816 bot815 bot816 {l}
Rtop_815_845 top815 top845 {r}
Ltop_815_845 top815 top845 {l}
Rbot_815_845 bot815 bot845 {r}
Lbot_815_845 bot815 bot845 {l}
C815 top815 bot815 {c}
Rtop_816_817 top816 top817 {r}
Ltop_816_817 top816 top817 {l}
Rbot_816_817 bot816 bot817 {r}
Lbot_816_817 bot816 bot817 {l}
Rtop_816_846 top816 top846 {r}
Ltop_816_846 top816 top846 {l}
Rbot_816_846 bot816 bot846 {r}
Lbot_816_846 bot816 bot846 {l}
C816 top816 bot816 {c}
Rtop_817_818 top817 top818 {r}
Ltop_817_818 top817 top818 {l}
Rbot_817_818 bot817 bot818 {r}
Lbot_817_818 bot817 bot818 {l}
Rtop_817_847 top817 top847 {r}
Ltop_817_847 top817 top847 {l}
Rbot_817_847 bot817 bot847 {r}
Lbot_817_847 bot817 bot847 {l}
C817 top817 bot817 {c}
Rtop_818_819 top818 top819 {r}
Ltop_818_819 top818 top819 {l}
Rbot_818_819 bot818 bot819 {r}
Lbot_818_819 bot818 bot819 {l}
Rtop_818_848 top818 top848 {r}
Ltop_818_848 top818 top848 {l}
Rbot_818_848 bot818 bot848 {r}
Lbot_818_848 bot818 bot848 {l}
C818 top818 bot818 {c}
Rtop_819_820 top819 top820 {r}
Ltop_819_820 top819 top820 {l}
Rbot_819_820 bot819 bot820 {r}
Lbot_819_820 bot819 bot820 {l}
Rtop_819_849 top819 top849 {r}
Ltop_819_849 top819 top849 {l}
Rbot_819_849 bot819 bot849 {r}
Lbot_819_849 bot819 bot849 {l}
C819 top819 bot819 {c}
Rtop_820_821 top820 top821 {r}
Ltop_820_821 top820 top821 {l}
Rbot_820_821 bot820 bot821 {r}
Lbot_820_821 bot820 bot821 {l}
Rtop_820_850 top820 top850 {r}
Ltop_820_850 top820 top850 {l}
Rbot_820_850 bot820 bot850 {r}
Lbot_820_850 bot820 bot850 {l}
C820 top820 bot820 {c}
Rtop_821_822 top821 top822 {r}
Ltop_821_822 top821 top822 {l}
Rbot_821_822 bot821 bot822 {r}
Lbot_821_822 bot821 bot822 {l}
Rtop_821_851 top821 top851 {r}
Ltop_821_851 top821 top851 {l}
Rbot_821_851 bot821 bot851 {r}
Lbot_821_851 bot821 bot851 {l}
C821 top821 bot821 {c}
Rtop_822_823 top822 top823 {r}
Ltop_822_823 top822 top823 {l}
Rbot_822_823 bot822 bot823 {r}
Lbot_822_823 bot822 bot823 {l}
Rtop_822_852 top822 top852 {r}
Ltop_822_852 top822 top852 {l}
Rbot_822_852 bot822 bot852 {r}
Lbot_822_852 bot822 bot852 {l}
C822 top822 bot822 {c}
Rtop_823_824 top823 top824 {r}
Ltop_823_824 top823 top824 {l}
Rbot_823_824 bot823 bot824 {r}
Lbot_823_824 bot823 bot824 {l}
Rtop_823_853 top823 top853 {r}
Ltop_823_853 top823 top853 {l}
Rbot_823_853 bot823 bot853 {r}
Lbot_823_853 bot823 bot853 {l}
C823 top823 bot823 {c}
Rtop_824_825 top824 top825 {r}
Ltop_824_825 top824 top825 {l}
Rbot_824_825 bot824 bot825 {r}
Lbot_824_825 bot824 bot825 {l}
Rtop_824_854 top824 top854 {r}
Ltop_824_854 top824 top854 {l}
Rbot_824_854 bot824 bot854 {r}
Lbot_824_854 bot824 bot854 {l}
C824 top824 bot824 {c}
Rtop_825_826 top825 top826 {r}
Ltop_825_826 top825 top826 {l}
Rbot_825_826 bot825 bot826 {r}
Lbot_825_826 bot825 bot826 {l}
Rtop_825_855 top825 top855 {r}
Ltop_825_855 top825 top855 {l}
Rbot_825_855 bot825 bot855 {r}
Lbot_825_855 bot825 bot855 {l}
C825 top825 bot825 {c}
Rtop_826_827 top826 top827 {r}
Ltop_826_827 top826 top827 {l}
Rbot_826_827 bot826 bot827 {r}
Lbot_826_827 bot826 bot827 {l}
Rtop_826_856 top826 top856 {r}
Ltop_826_856 top826 top856 {l}
Rbot_826_856 bot826 bot856 {r}
Lbot_826_856 bot826 bot856 {l}
C826 top826 bot826 {c}
Rtop_827_828 top827 top828 {r}
Ltop_827_828 top827 top828 {l}
Rbot_827_828 bot827 bot828 {r}
Lbot_827_828 bot827 bot828 {l}
Rtop_827_857 top827 top857 {r}
Ltop_827_857 top827 top857 {l}
Rbot_827_857 bot827 bot857 {r}
Lbot_827_857 bot827 bot857 {l}
C827 top827 bot827 {c}
Rtop_828_829 top828 top829 {r}
Ltop_828_829 top828 top829 {l}
Rbot_828_829 bot828 bot829 {r}
Lbot_828_829 bot828 bot829 {l}
Rtop_828_858 top828 top858 {r}
Ltop_828_858 top828 top858 {l}
Rbot_828_858 bot828 bot858 {r}
Lbot_828_858 bot828 bot858 {l}
C828 top828 bot828 {c}
Rtop_829_830 top829 top830 {r}
Ltop_829_830 top829 top830 {l}
Rbot_829_830 bot829 bot830 {r}
Lbot_829_830 bot829 bot830 {l}
Rtop_829_859 top829 top859 {r}
Ltop_829_859 top829 top859 {l}
Rbot_829_859 bot829 bot859 {r}
Lbot_829_859 bot829 bot859 {l}
C829 top829 bot829 {c}
Rtop_830_831 top830 top831 {r}
Ltop_830_831 top830 top831 {l}
Rbot_830_831 bot830 bot831 {r}
Lbot_830_831 bot830 bot831 {l}
Rtop_830_860 top830 top860 {r}
Ltop_830_860 top830 top860 {l}
Rbot_830_860 bot830 bot860 {r}
Lbot_830_860 bot830 bot860 {l}
C830 top830 bot830 {c}
Rtop_831_832 top831 top832 {r}
Ltop_831_832 top831 top832 {l}
Rbot_831_832 bot831 bot832 {r}
Lbot_831_832 bot831 bot832 {l}
Rtop_831_861 top831 top861 {r}
Ltop_831_861 top831 top861 {l}
Rbot_831_861 bot831 bot861 {r}
Lbot_831_861 bot831 bot861 {l}
C831 top831 bot831 {c}
Rtop_832_833 top832 top833 {r}
Ltop_832_833 top832 top833 {l}
Rbot_832_833 bot832 bot833 {r}
Lbot_832_833 bot832 bot833 {l}
Rtop_832_862 top832 top862 {r}
Ltop_832_862 top832 top862 {l}
Rbot_832_862 bot832 bot862 {r}
Lbot_832_862 bot832 bot862 {l}
C832 top832 bot832 {c}
Rtop_833_834 top833 top834 {r}
Ltop_833_834 top833 top834 {l}
Rbot_833_834 bot833 bot834 {r}
Lbot_833_834 bot833 bot834 {l}
Rtop_833_863 top833 top863 {r}
Ltop_833_863 top833 top863 {l}
Rbot_833_863 bot833 bot863 {r}
Lbot_833_863 bot833 bot863 {l}
C833 top833 bot833 {c}
Rtop_834_835 top834 top835 {r}
Ltop_834_835 top834 top835 {l}
Rbot_834_835 bot834 bot835 {r}
Lbot_834_835 bot834 bot835 {l}
Rtop_834_864 top834 top864 {r}
Ltop_834_864 top834 top864 {l}
Rbot_834_864 bot834 bot864 {r}
Lbot_834_864 bot834 bot864 {l}
C834 top834 bot834 {c}
Rtop_835_836 top835 top836 {r}
Ltop_835_836 top835 top836 {l}
Rbot_835_836 bot835 bot836 {r}
Lbot_835_836 bot835 bot836 {l}
Rtop_835_865 top835 top865 {r}
Ltop_835_865 top835 top865 {l}
Rbot_835_865 bot835 bot865 {r}
Lbot_835_865 bot835 bot865 {l}
C835 top835 bot835 {c}
Rtop_836_837 top836 top837 {r}
Ltop_836_837 top836 top837 {l}
Rbot_836_837 bot836 bot837 {r}
Lbot_836_837 bot836 bot837 {l}
Rtop_836_866 top836 top866 {r}
Ltop_836_866 top836 top866 {l}
Rbot_836_866 bot836 bot866 {r}
Lbot_836_866 bot836 bot866 {l}
C836 top836 bot836 {c}
Rtop_837_838 top837 top838 {r}
Ltop_837_838 top837 top838 {l}
Rbot_837_838 bot837 bot838 {r}
Lbot_837_838 bot837 bot838 {l}
Rtop_837_867 top837 top867 {r}
Ltop_837_867 top837 top867 {l}
Rbot_837_867 bot837 bot867 {r}
Lbot_837_867 bot837 bot867 {l}
C837 top837 bot837 {c}
Rtop_838_839 top838 top839 {r}
Ltop_838_839 top838 top839 {l}
Rbot_838_839 bot838 bot839 {r}
Lbot_838_839 bot838 bot839 {l}
Rtop_838_868 top838 top868 {r}
Ltop_838_868 top838 top868 {l}
Rbot_838_868 bot838 bot868 {r}
Lbot_838_868 bot838 bot868 {l}
C838 top838 bot838 {c}
Rtop_839_840 top839 top840 {r}
Ltop_839_840 top839 top840 {l}
Rbot_839_840 bot839 bot840 {r}
Lbot_839_840 bot839 bot840 {l}
Rtop_839_869 top839 top869 {r}
Ltop_839_869 top839 top869 {l}
Rbot_839_869 bot839 bot869 {r}
Lbot_839_869 bot839 bot869 {l}
C839 top839 bot839 {c}
Rtop_840_870 top840 top870 {r}
Ltop_840_870 top840 top870 {l}
Rbot_840_870 bot840 bot870 {r}
Lbot_840_870 bot840 bot870 {l}
C840 top840 bot840 {c}
Rtop_841_842 top841 top842 {r}
Ltop_841_842 top841 top842 {l}
Rbot_841_842 bot841 bot842 {r}
Lbot_841_842 bot841 bot842 {l}
Rtop_841_871 top841 top871 {r}
Ltop_841_871 top841 top871 {l}
Rbot_841_871 bot841 bot871 {r}
Lbot_841_871 bot841 bot871 {l}
C841 top841 bot841 {c}
Rtop_842_843 top842 top843 {r}
Ltop_842_843 top842 top843 {l}
Rbot_842_843 bot842 bot843 {r}
Lbot_842_843 bot842 bot843 {l}
Rtop_842_872 top842 top872 {r}
Ltop_842_872 top842 top872 {l}
Rbot_842_872 bot842 bot872 {r}
Lbot_842_872 bot842 bot872 {l}
C842 top842 bot842 {c}
Rtop_843_844 top843 top844 {r}
Ltop_843_844 top843 top844 {l}
Rbot_843_844 bot843 bot844 {r}
Lbot_843_844 bot843 bot844 {l}
Rtop_843_873 top843 top873 {r}
Ltop_843_873 top843 top873 {l}
Rbot_843_873 bot843 bot873 {r}
Lbot_843_873 bot843 bot873 {l}
C843 top843 bot843 {c}
Rtop_844_845 top844 top845 {r}
Ltop_844_845 top844 top845 {l}
Rbot_844_845 bot844 bot845 {r}
Lbot_844_845 bot844 bot845 {l}
Rtop_844_874 top844 top874 {r}
Ltop_844_874 top844 top874 {l}
Rbot_844_874 bot844 bot874 {r}
Lbot_844_874 bot844 bot874 {l}
C844 top844 bot844 {c}
Rtop_845_846 top845 top846 {r}
Ltop_845_846 top845 top846 {l}
Rbot_845_846 bot845 bot846 {r}
Lbot_845_846 bot845 bot846 {l}
Rtop_845_875 top845 top875 {r}
Ltop_845_875 top845 top875 {l}
Rbot_845_875 bot845 bot875 {r}
Lbot_845_875 bot845 bot875 {l}
C845 top845 bot845 {c}
Rtop_846_847 top846 top847 {r}
Ltop_846_847 top846 top847 {l}
Rbot_846_847 bot846 bot847 {r}
Lbot_846_847 bot846 bot847 {l}
Rtop_846_876 top846 top876 {r}
Ltop_846_876 top846 top876 {l}
Rbot_846_876 bot846 bot876 {r}
Lbot_846_876 bot846 bot876 {l}
C846 top846 bot846 {c}
Rtop_847_848 top847 top848 {r}
Ltop_847_848 top847 top848 {l}
Rbot_847_848 bot847 bot848 {r}
Lbot_847_848 bot847 bot848 {l}
Rtop_847_877 top847 top877 {r}
Ltop_847_877 top847 top877 {l}
Rbot_847_877 bot847 bot877 {r}
Lbot_847_877 bot847 bot877 {l}
C847 top847 bot847 {c}
Rtop_848_849 top848 top849 {r}
Ltop_848_849 top848 top849 {l}
Rbot_848_849 bot848 bot849 {r}
Lbot_848_849 bot848 bot849 {l}
Rtop_848_878 top848 top878 {r}
Ltop_848_878 top848 top878 {l}
Rbot_848_878 bot848 bot878 {r}
Lbot_848_878 bot848 bot878 {l}
C848 top848 bot848 {c}
Rtop_849_850 top849 top850 {r}
Ltop_849_850 top849 top850 {l}
Rbot_849_850 bot849 bot850 {r}
Lbot_849_850 bot849 bot850 {l}
Rtop_849_879 top849 top879 {r}
Ltop_849_879 top849 top879 {l}
Rbot_849_879 bot849 bot879 {r}
Lbot_849_879 bot849 bot879 {l}
C849 top849 bot849 {c}
Rtop_850_851 top850 top851 {r}
Ltop_850_851 top850 top851 {l}
Rbot_850_851 bot850 bot851 {r}
Lbot_850_851 bot850 bot851 {l}
Rtop_850_880 top850 top880 {r}
Ltop_850_880 top850 top880 {l}
Rbot_850_880 bot850 bot880 {r}
Lbot_850_880 bot850 bot880 {l}
C850 top850 bot850 {c}
Rtop_851_852 top851 top852 {r}
Ltop_851_852 top851 top852 {l}
Rbot_851_852 bot851 bot852 {r}
Lbot_851_852 bot851 bot852 {l}
Rtop_851_881 top851 top881 {r}
Ltop_851_881 top851 top881 {l}
Rbot_851_881 bot851 bot881 {r}
Lbot_851_881 bot851 bot881 {l}
C851 top851 bot851 {c}
Rtop_852_853 top852 top853 {r}
Ltop_852_853 top852 top853 {l}
Rbot_852_853 bot852 bot853 {r}
Lbot_852_853 bot852 bot853 {l}
Rtop_852_882 top852 top882 {r}
Ltop_852_882 top852 top882 {l}
Rbot_852_882 bot852 bot882 {r}
Lbot_852_882 bot852 bot882 {l}
C852 top852 bot852 {c}
Rtop_853_854 top853 top854 {r}
Ltop_853_854 top853 top854 {l}
Rbot_853_854 bot853 bot854 {r}
Lbot_853_854 bot853 bot854 {l}
Rtop_853_883 top853 top883 {r}
Ltop_853_883 top853 top883 {l}
Rbot_853_883 bot853 bot883 {r}
Lbot_853_883 bot853 bot883 {l}
C853 top853 bot853 {c}
Rtop_854_855 top854 top855 {r}
Ltop_854_855 top854 top855 {l}
Rbot_854_855 bot854 bot855 {r}
Lbot_854_855 bot854 bot855 {l}
Rtop_854_884 top854 top884 {r}
Ltop_854_884 top854 top884 {l}
Rbot_854_884 bot854 bot884 {r}
Lbot_854_884 bot854 bot884 {l}
C854 top854 bot854 {c}
Rtop_855_856 top855 top856 {r}
Ltop_855_856 top855 top856 {l}
Rbot_855_856 bot855 bot856 {r}
Lbot_855_856 bot855 bot856 {l}
Rtop_855_885 top855 top885 {r}
Ltop_855_885 top855 top885 {l}
Rbot_855_885 bot855 bot885 {r}
Lbot_855_885 bot855 bot885 {l}
C855 top855 bot855 {c}
Rtop_856_857 top856 top857 {r}
Ltop_856_857 top856 top857 {l}
Rbot_856_857 bot856 bot857 {r}
Lbot_856_857 bot856 bot857 {l}
Rtop_856_886 top856 top886 {r}
Ltop_856_886 top856 top886 {l}
Rbot_856_886 bot856 bot886 {r}
Lbot_856_886 bot856 bot886 {l}
C856 top856 bot856 {c}
Rtop_857_858 top857 top858 {r}
Ltop_857_858 top857 top858 {l}
Rbot_857_858 bot857 bot858 {r}
Lbot_857_858 bot857 bot858 {l}
Rtop_857_887 top857 top887 {r}
Ltop_857_887 top857 top887 {l}
Rbot_857_887 bot857 bot887 {r}
Lbot_857_887 bot857 bot887 {l}
C857 top857 bot857 {c}
Rtop_858_859 top858 top859 {r}
Ltop_858_859 top858 top859 {l}
Rbot_858_859 bot858 bot859 {r}
Lbot_858_859 bot858 bot859 {l}
Rtop_858_888 top858 top888 {r}
Ltop_858_888 top858 top888 {l}
Rbot_858_888 bot858 bot888 {r}
Lbot_858_888 bot858 bot888 {l}
C858 top858 bot858 {c}
Rtop_859_860 top859 top860 {r}
Ltop_859_860 top859 top860 {l}
Rbot_859_860 bot859 bot860 {r}
Lbot_859_860 bot859 bot860 {l}
Rtop_859_889 top859 top889 {r}
Ltop_859_889 top859 top889 {l}
Rbot_859_889 bot859 bot889 {r}
Lbot_859_889 bot859 bot889 {l}
C859 top859 bot859 {c}
Rtop_860_861 top860 top861 {r}
Ltop_860_861 top860 top861 {l}
Rbot_860_861 bot860 bot861 {r}
Lbot_860_861 bot860 bot861 {l}
Rtop_860_890 top860 top890 {r}
Ltop_860_890 top860 top890 {l}
Rbot_860_890 bot860 bot890 {r}
Lbot_860_890 bot860 bot890 {l}
C860 top860 bot860 {c}
Rtop_861_862 top861 top862 {r}
Ltop_861_862 top861 top862 {l}
Rbot_861_862 bot861 bot862 {r}
Lbot_861_862 bot861 bot862 {l}
Rtop_861_891 top861 top891 {r}
Ltop_861_891 top861 top891 {l}
Rbot_861_891 bot861 bot891 {r}
Lbot_861_891 bot861 bot891 {l}
C861 top861 bot861 {c}
Rtop_862_863 top862 top863 {r}
Ltop_862_863 top862 top863 {l}
Rbot_862_863 bot862 bot863 {r}
Lbot_862_863 bot862 bot863 {l}
Rtop_862_892 top862 top892 {r}
Ltop_862_892 top862 top892 {l}
Rbot_862_892 bot862 bot892 {r}
Lbot_862_892 bot862 bot892 {l}
C862 top862 bot862 {c}
Rtop_863_864 top863 top864 {r}
Ltop_863_864 top863 top864 {l}
Rbot_863_864 bot863 bot864 {r}
Lbot_863_864 bot863 bot864 {l}
Rtop_863_893 top863 top893 {r}
Ltop_863_893 top863 top893 {l}
Rbot_863_893 bot863 bot893 {r}
Lbot_863_893 bot863 bot893 {l}
C863 top863 bot863 {c}
Rtop_864_865 top864 top865 {r}
Ltop_864_865 top864 top865 {l}
Rbot_864_865 bot864 bot865 {r}
Lbot_864_865 bot864 bot865 {l}
Rtop_864_894 top864 top894 {r}
Ltop_864_894 top864 top894 {l}
Rbot_864_894 bot864 bot894 {r}
Lbot_864_894 bot864 bot894 {l}
C864 top864 bot864 {c}
Rtop_865_866 top865 top866 {r}
Ltop_865_866 top865 top866 {l}
Rbot_865_866 bot865 bot866 {r}
Lbot_865_866 bot865 bot866 {l}
Rtop_865_895 top865 top895 {r}
Ltop_865_895 top865 top895 {l}
Rbot_865_895 bot865 bot895 {r}
Lbot_865_895 bot865 bot895 {l}
C865 top865 bot865 {c}
Rtop_866_867 top866 top867 {r}
Ltop_866_867 top866 top867 {l}
Rbot_866_867 bot866 bot867 {r}
Lbot_866_867 bot866 bot867 {l}
Rtop_866_896 top866 top896 {r}
Ltop_866_896 top866 top896 {l}
Rbot_866_896 bot866 bot896 {r}
Lbot_866_896 bot866 bot896 {l}
C866 top866 bot866 {c}
Rtop_867_868 top867 top868 {r}
Ltop_867_868 top867 top868 {l}
Rbot_867_868 bot867 bot868 {r}
Lbot_867_868 bot867 bot868 {l}
Rtop_867_897 top867 top897 {r}
Ltop_867_897 top867 top897 {l}
Rbot_867_897 bot867 bot897 {r}
Lbot_867_897 bot867 bot897 {l}
C867 top867 bot867 {c}
Rtop_868_869 top868 top869 {r}
Ltop_868_869 top868 top869 {l}
Rbot_868_869 bot868 bot869 {r}
Lbot_868_869 bot868 bot869 {l}
Rtop_868_898 top868 top898 {r}
Ltop_868_898 top868 top898 {l}
Rbot_868_898 bot868 bot898 {r}
Lbot_868_898 bot868 bot898 {l}
C868 top868 bot868 {c}
Rtop_869_870 top869 top870 {r}
Ltop_869_870 top869 top870 {l}
Rbot_869_870 bot869 bot870 {r}
Lbot_869_870 bot869 bot870 {l}
Rtop_869_899 top869 top899 {r}
Ltop_869_899 top869 top899 {l}
Rbot_869_899 bot869 bot899 {r}
Lbot_869_899 bot869 bot899 {l}
C869 top869 bot869 {c}
Rtop_870_900 top870 top900 {r}
Ltop_870_900 top870 top900 {l}
Rbot_870_900 bot870 bot900 {r}
Lbot_870_900 bot870 bot900 {l}
C870 top870 bot870 {c}
Rtop_871_872 top871 top872 {r}
Ltop_871_872 top871 top872 {l}
Rbot_871_872 bot871 bot872 {r}
Lbot_871_872 bot871 bot872 {l}
C871 top871 bot871 {c}
Rtop_872_873 top872 top873 {r}
Ltop_872_873 top872 top873 {l}
Rbot_872_873 bot872 bot873 {r}
Lbot_872_873 bot872 bot873 {l}
C872 top872 bot872 {c}
Rtop_873_874 top873 top874 {r}
Ltop_873_874 top873 top874 {l}
Rbot_873_874 bot873 bot874 {r}
Lbot_873_874 bot873 bot874 {l}
C873 top873 bot873 {c}
Rtop_874_875 top874 top875 {r}
Ltop_874_875 top874 top875 {l}
Rbot_874_875 bot874 bot875 {r}
Lbot_874_875 bot874 bot875 {l}
C874 top874 bot874 {c}
Rtop_875_876 top875 top876 {r}
Ltop_875_876 top875 top876 {l}
Rbot_875_876 bot875 bot876 {r}
Lbot_875_876 bot875 bot876 {l}
C875 top875 bot875 {c}
Rtop_876_877 top876 top877 {r}
Ltop_876_877 top876 top877 {l}
Rbot_876_877 bot876 bot877 {r}
Lbot_876_877 bot876 bot877 {l}
C876 top876 bot876 {c}
Rtop_877_878 top877 top878 {r}
Ltop_877_878 top877 top878 {l}
Rbot_877_878 bot877 bot878 {r}
Lbot_877_878 bot877 bot878 {l}
C877 top877 bot877 {c}
Rtop_878_879 top878 top879 {r}
Ltop_878_879 top878 top879 {l}
Rbot_878_879 bot878 bot879 {r}
Lbot_878_879 bot878 bot879 {l}
C878 top878 bot878 {c}
Rtop_879_880 top879 top880 {r}
Ltop_879_880 top879 top880 {l}
Rbot_879_880 bot879 bot880 {r}
Lbot_879_880 bot879 bot880 {l}
C879 top879 bot879 {c}
Rtop_880_881 top880 top881 {r}
Ltop_880_881 top880 top881 {l}
Rbot_880_881 bot880 bot881 {r}
Lbot_880_881 bot880 bot881 {l}
C880 top880 bot880 {c}
Rtop_881_882 top881 top882 {r}
Ltop_881_882 top881 top882 {l}
Rbot_881_882 bot881 bot882 {r}
Lbot_881_882 bot881 bot882 {l}
C881 top881 bot881 {c}
Rtop_882_883 top882 top883 {r}
Ltop_882_883 top882 top883 {l}
Rbot_882_883 bot882 bot883 {r}
Lbot_882_883 bot882 bot883 {l}
C882 top882 bot882 {c}
Rtop_883_884 top883 top884 {r}
Ltop_883_884 top883 top884 {l}
Rbot_883_884 bot883 bot884 {r}
Lbot_883_884 bot883 bot884 {l}
C883 top883 bot883 {c}
Rtop_884_885 top884 top885 {r}
Ltop_884_885 top884 top885 {l}
Rbot_884_885 bot884 bot885 {r}
Lbot_884_885 bot884 bot885 {l}
C884 top884 bot884 {c}
Rtop_885_886 top885 top886 {r}
Ltop_885_886 top885 top886 {l}
Rbot_885_886 bot885 bot886 {r}
Lbot_885_886 bot885 bot886 {l}
C885 top885 bot885 {c}
Rtop_886_887 top886 top887 {r}
Ltop_886_887 top886 top887 {l}
Rbot_886_887 bot886 bot887 {r}
Lbot_886_887 bot886 bot887 {l}
C886 top886 bot886 {c}
Rtop_887_888 top887 top888 {r}
Ltop_887_888 top887 top888 {l}
Rbot_887_888 bot887 bot888 {r}
Lbot_887_888 bot887 bot888 {l}
C887 top887 bot887 {c}
Rtop_888_889 top888 top889 {r}
Ltop_888_889 top888 top889 {l}
Rbot_888_889 bot888 bot889 {r}
Lbot_888_889 bot888 bot889 {l}
C888 top888 bot888 {c}
Rtop_889_890 top889 top890 {r}
Ltop_889_890 top889 top890 {l}
Rbot_889_890 bot889 bot890 {r}
Lbot_889_890 bot889 bot890 {l}
C889 top889 bot889 {c}
Rtop_890_891 top890 top891 {r}
Ltop_890_891 top890 top891 {l}
Rbot_890_891 bot890 bot891 {r}
Lbot_890_891 bot890 bot891 {l}
C890 top890 bot890 {c}
Rtop_891_892 top891 top892 {r}
Ltop_891_892 top891 top892 {l}
Rbot_891_892 bot891 bot892 {r}
Lbot_891_892 bot891 bot892 {l}
C891 top891 bot891 {c}
Rtop_892_893 top892 top893 {r}
Ltop_892_893 top892 top893 {l}
Rbot_892_893 bot892 bot893 {r}
Lbot_892_893 bot892 bot893 {l}
C892 top892 bot892 {c}
Rtop_893_894 top893 top894 {r}
Ltop_893_894 top893 top894 {l}
Rbot_893_894 bot893 bot894 {r}
Lbot_893_894 bot893 bot894 {l}
C893 top893 bot893 {c}
Rtop_894_895 top894 top895 {r}
Ltop_894_895 top894 top895 {l}
Rbot_894_895 bot894 bot895 {r}
Lbot_894_895 bot894 bot895 {l}
C894 top894 bot894 {c}
Rtop_895_896 top895 top896 {r}
Ltop_895_896 top895 top896 {l}
Rbot_895_896 bot895 bot896 {r}
Lbot_895_896 bot895 bot896 {l}
C895 top895 bot895 {c}
Rtop_896_897 top896 top897 {r}
Ltop_896_897 top896 top897 {l}
Rbot_896_897 bot896 bot897 {r}
Lbot_896_897 bot896 bot897 {l}
C896 top896 bot896 {c}
Rtop_897_898 top897 top898 {r}
Ltop_897_898 top897 top898 {l}
Rbot_897_898 bot897 bot898 {r}
Lbot_897_898 bot897 bot898 {l}
C897 top897 bot897 {c}
Rtop_898_899 top898 top899 {r}
Ltop_898_899 top898 top899 {l}
Rbot_898_899 bot898 bot899 {r}
Lbot_898_899 bot898 bot899 {l}
C898 top898 bot898 {c}
Rtop_899_900 top899 top900 {r}
Ltop_899_900 top899 top900 {l}
Rbot_899_900 bot899 bot900 {r}
Lbot_899_900 bot899 bot900 {l}
C899 top899 bot899 {c}
C900 top900 bot900 {c}
.ends

X1 in out 0 grids
v1 in 0 ac 1 dc 0

*>.print ac vr(out) vi(out) vm(out) vp(out)
*>.print op v(out)
*>.op
*>.ac oct 1 1 250k basic
*>.status notime
*>.end

* try this with ngspice -b ..
.control
ac oct 1 1 500k
set units = degrees
.endc
.print ac vm(out) vp(out)
