
.model foo d
x1 (a b c) foo
.op
.end
