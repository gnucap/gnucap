# PWL sources
v1 1 0 PWL  0,0 1,1 4,2 9,3 16,4 25,5
i1 2 0 PWL  0,0 1,-1 4,2 9,-3 16,4 25,-5
r4 2 0 10k
.list
.print op v(nodes)
.op
.print dc v(nodes)
.dc v1 -10 10 1
.print tran v(nodes)
.tran 0 30 1
.end
