* int vs float check
.param  x='3+a+1.+1'
.eval x
.eval 3.+a+1+1
.eval a+b
.eval 2+a+b+3
.eval a+2+b+3
.eval a+2+3+b
.eval 2+a+3+b
.eval 2/a
.eval 2/3
.eval 2/3.
.eval 2./3
.param a=2.
.eval x
.eval 3+a+1+1
.eval a+b
.eval 2+a+b+3
.eval a+2+b+3
.eval a+2+3+b
.eval 2+a+3+b
.eval a/3
.param a=3
.eval a
.eval 3/3
.eval a/3
.eval 0 + 0.
.eval 0 + 0
.eval 4 + 0.
.eval 1/2
.eval (-5)/2
.end
