'inductance check, no tolerance
V1   1  0  dc 1 ac 1
L3   1  2  1.
R4   2  0  1.
R5   1  3  1.
C6   3  0  1.
.print dc v(3)
.print ac v(3)
.dc v1 1 10 1
.ac dec 10 .1 10
.status notime
.end
