A 9217 node circuit
Vin 1 0 dc sin 0 1 1k 0 0
x1 1 2 eq64
x2 2 3 eq64
x3 3 4 eq64
x4 4 5 eq64
.subckt eq64 1 5
x1 1 2 eq16
x2 2 3 eq16
x3 3 4 eq16
x4 4 5 eq16
.ends eq64
.subckt eq16 1 5
x1 1 2 eq4
x2 2 3 eq4
x3 3 4 eq4
x4 4 5 eq4
.ends eq16
.subckt eq4 1 5
x1 1 2 eq
x2 2 3 eq
x3 3 4 eq
x4 4 5 eq
.ends eq4
.subckt eq 31 37
R101a   35   1  50.K
R101b   36   1  50.K
R102a   32   4  50.K
R102b   33   4  50.K
R103a   35   7  50.K
R103b   36   7  50.K
R104a   32  10  50.K
R104b   33  10  50.K
R105a   35  13  50.K
R105b   36  13  50.K
R106a   32  16  50.K
R106b   33  16  50.K
R107a   35  19  50.K
R107b   36  19  50.K
R108a   32  22  50.K
R108b   33  22  50.K
R109a   35  25  50.K
R109b   36  25  50.K
R110a   32  28  50.K
R110b   33  28  50.K
C1      1   2  1.5u
C2      4   5  748.n
C3      7   8  408.n
C4     10  11  206.n
C5     13  14  100.n
C6     16  17  50.9n
C7     19  20  25.3n
C8     22  23  12.7n
C9     25  26  5.9n
C10    28  29  2.95n
C11     2   3  15.n
C12     5   6  6.8n
C13     8   9  3.3n
C14    11  12  1.8n
C15    14  15  1.n
C16    17  18  470.p
C17    20  21  220.p
C18    23  24  120.p
C19    26  27  68.p
C20    29  30  33.p
R1      3   0  475.K
R2      6   0  536.K
R3      9   0  549.K
R4     12   0  499.K
R5     15   0  464.K
R6     18   0  475.K
R7     21   0  523.K
R8     24   0  475.K
R9     27   0  412.K
R10    30   0  422.K
G5a     2   0   3   0   -.000416666
R11     2   0  2.4K
G5b     5   0   6   0   -.000416666
R12     5   0  2.4K
G6a     8   0   9   0   -.000454545
R13     8   0  2.2K
G6b    11   0  12   0   -.000454545
R14    11   0  2.2K
G7a    14   0  15   0   -.000454545
R15    14   0  2.2K
G7b    17   0  18   0   -.000454545
R16    17   0  2.2K
G8a    20   0  21   0   -.000454545
R17    20   0  2.2K
G8b    23   0  24   0   -.000454545
R18    23   0  2.2K
G9a    26   0  27   0   -.000416666
R19    26   0  2.4K
G9b    29   0  30   0   -.000416666
R20    29   0  2.4K
R29    31  32  9.1K
R30    33  34  9.1K
R31    34  35  9.1K
R32    36  37  9.1K
C25    31  32  150.p
C26    33  34  150.p
C27    34  35  150.p
C28    36  37  150.p
E2     34   0  32  33  10.K
E3     37   0  35  36  10.K
.option acct
.ends eq
.print tran v(5)
.tran .00001 .001 0 
.end
