
m1 3 2 0 0 foo
.model foo d
.op
.end
