bug, some models don't complain when parameters move out of range

.model nmos.1 nmos level=1 vto=0.7 lmin=1e-6 lmax=2e-6

Mn1 3 2 0 0 NMOS W=8e-6 L=L

.parameter L=1e-6
.dc
.parameter L=5e-6
.dc
.dc L 1e-6 3e-6 1e-6

.end
