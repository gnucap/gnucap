
.subckt foo (1 2)
r1 (1 2) 1
.ends
v1 (1 0) 1
x1 (1 2) foo
x2 (2 3) x1
.op
.list
.end
