'inductance check, no tolerance
V1   1  0  generator(1)
L3   1  2  1.
R4   2  0  1.
R5   1  3  .97
C6   3  0  1.
.options short=1p
.width out=170
.list
.print tran iter(0)  v(nodes) z(c6) zraw(c6) z(3)
.fanout
.fanout 2
.tran 0 1 .1
.print ac v(2) v(3) vp(2) vp(3) z(c6) zraw(c6) z(3)
.ac .001 10 decade 2
.list
.end
