' exp test, periodic
.option out=170
.param p=20n
v1 1 0 exp  iv= 0.  pv= 1.  td1=p/20  tau1=p/4  td2=p/2  tau2=p/4  period=p
.print tran v(1) next(v1) event(v1) control(0)
.tran 0 100n 100n trace all
.list
.end
