nonlinear res test

V1 1 0  1.
R1 1 0 PWL
+-102400,-1.1
+ -51200,-1.0
+ -25600, -.9
+ -12800, -.8
+  -6400, -.7
+  -3200, -.6
+  -1600, -.5
+   -800, -.4
+   -400, -.3
+   -200, -.2
+   -100, -.1
+  -.500, -.05
+      0,  .0
+   .500,  .05
+    100,  .1
+    200,  .2
+    400,  .3
+    800,  .4
+   1600,  .5
+   3200,  .6
+   6400,  .7
+  12800,  .8
+  25600,  .9
+  51200, 1.0
+102400, 1.1

*.options nopicky
.options short 1e-5
.print dc i(R1) vin(r1) i(v1) iter(0) f(R1) df(R1) in(R1) iof(R1)
.dc v1 -1 1 0.1 loop trace n basic > res.out
.stat notime
