' test nested subckts
.option trace
.subckt aa (a b c)
.subckt bb (1 2)
r1 (1 2) 1k
.ends bb
r1 (a b) 1
r2 (b 0) 1
r3 (b c) 1
xh (a b) bb
.ends aa
x1 (1 2 3) aa
v1 (1 0) dc 1
.list
.print op v(nodes)
.op
.end
