
v1 2 0 sin freq=1k
d1 0 2 dd
w3 1 0 d1 foo
r3 1 3 1k
v3 3 0 dc 1
.model foo csw
.model dd d
.probe tran v(nodes) iter(0)
.tran 0 .002 100u
.end
