TRANSFER curve tracer, ig-spice
*
* Sources that we sweep
VIN 1 0 1
*VOUT 2 0 5
VBACK 0 6 0
EBACK 7 5 0 6 1
*
* power supplies, etc.
VDD 5 0 5
*
* "ammeters" (fudge)
*VPU 3 2 0
*VPD 2 4 0
VPU 3 0 0
VPD 5 4 0
*
* active devices
MPU 3 1 5 7 CMOSP L=3U W=6U AD=18P AS=18P PD=18U PS=18U
MPD 4 1 0 6 CMOSN L=3U W=3U AD=9P AS=9P PD=12U PS=12U
*
* models
.MODEL CMOSN NMOS LEVEL=2 LD=0.265073U TOX=418.0E-10
+ NSUB=1.53142E+16 VTO=0.844345 KP=4.15964E-05 GAMMA=0.863074
+ PHI=0.6 UO=503.521 UEXP=0.163917 UCRIT=161166
+ DELTA=1E-06 VMAX=55903.5 XJ=0.400000U LAMBDA=0.00906241
+ NFS=3.5934E+12 NEFF=1.001 NSS=1E+12 TPG=1.000000
+ RSH=0 CGDO=2.18971E-10 CGSO=2.18971E-10
+ CJ=0.0003844 MJ=0.488400 CJSW=5.272E-10 MJSW=0.300200 PB=0.700000
*
.MODEL CMOSP PMOS LEVEL=2 LD=0.299878U TOX=418.0E-10
+ NSUB=4.19363E+15 VTO=-0.79089 KP=1.64047E-05 GAMMA=0.451645
+ PHI=0.6 UO=198.577 UEXP=0.343935 UCRIT=110988
+ DELTA=0.956806 VMAX=41456.3 XJ=0.400000U LAMBDA=0.0344407
+ NFS=1E+12 NEFF=1.001 NSS=1E+12 TPG=-1.000000
+ RSH=0 CGDO=2.47722E-10 CGSO=2.47722E-10
+ CJ=0.0002281 MJ=0.508000 CJSW=3.077E-10 MJSW=0.193500 PB=0.740000
*
.OPTIONS LIMPTS=1000
.print op V(1) V(6) I(VPU) I(VPD) id(MPU) id(MPD) iter(0)
.print DC V(1) V(6) I(VPU) I(VPD) id(MPU) id(MPD) iter(0)
.op
.DC VDD 0 5 1 VIN 0 5 1
.DC VIN 0 5 1 VBACK 0 5 1
*>.status notime
.END
