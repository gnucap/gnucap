'nothing
.status
.end
