' test file for ap_ctof.cc
V1 1 0 1
R0102 1 2 -21.33t
R0200 2 0 7.3g
R0203 2 3 2.3k
R0300 3 0 3.4f
R0304 3 4 -3.4443323223p
R0400 4 0 4534445.3n
R0405 4 5 .23423u
R0500 5 0 -.000000000004343m
R0506 5 6 345345345Meg
R0600 6 0 23.432mil
R0607 6 7 4.55e-3
R0700 7 0 -344e28
R0708 7 8 0000004737e+77
R0800 8 0 -344e+28
R0809 8 9 +344e+28
R0900 9 0 foo
.list
.end
