# cccs test
i1 1 0 dc 11 ac 11
ri1 1 0 10
e1 2 0 1 0 8
re1 2 0 10
# sense the voltage source (0 volts)
i2 3 0 dc 11 ac 11
ri2 4 0 10
v2 3 4 0
h2 5 0 v2 8
rh2 5 0 10
# sense the resistor
i3 6 0 dc 11 ac 11
ri3 7 0 10
v3 6 7 0
h3 8 0 ri3 8
rh3 8 0 10
# sense the current source
i4 9 0 dc 11 ac 11
ri4 10 0 10
v4 9 10 0
h4 11 0 i4 8
rh4 11 0 10
# sense a conductance
i5 12 0 dc 11 ac 11
yi5 13 0 10
v5 12 13 0
h5 14 0 yi5 8
rh5 14 0 10
# sense a vccs
v6 15 0 dc 1.1 ac 1.1
g6 16 0 15 0 10
yi6 17 0 10
v6 16 17 0
h6 18 0 yi6 8
rh6 18 0 10
# sense a live voltage source
v7 19 0 dc 11 ac 11
rv7 19 0 10
h7 20 0 v7 8
rh7 20 0 10
# sense the resistor in series
v8 21 0 dc 11 ac 11
rv8 21 0 10
h8 22 0 rv8 8
rh8 22 0 10
# sense a vcvs
v9 23 0 dc 1.1 ac 1.1
e9 24 0 23 0 10
re9 24 0 10
h9a 25 0 e9 10
rh9a 25 0 10
h9b 26 0 re9 10
rh9b 26 0 10

.opt out 160
.print op v(nodes) i(v7) i(v8) i(e9) i(re9)
.op
.print tran v(nodes) i(v7) i(v8) i(e9) i(re9)
.tran 0 .1 .05
.print ac v(nodes) i(v7) i(v8) i(e9) i(re9)
.ac 1k
.end
