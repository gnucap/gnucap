'hyperbolic tangent test circuit
v1 1 0 generator(1)
e1 2 0 1 0 tanh 5 5
e2 3 0 1 0 tanh gain -5 limit 3
e3 4 0 1 0 tanh 4 limit 3
.print dc v nodes
.print ac v nodes
.dc -2 2 .1
.ac
.dc 1
.ac
.dc 0
.ac
.dc 1000
.ac
.list
.end
