'lib test

.lib test1
r1 (1 2) 1
.endl test1

.lib test2
v1 (1 0) 1
.lib c_lib.1.ckt test1
r2 (2 0) 1
.endl

r3 (2 3) 10k
r4 (3 0) 10k
.lib c_lib.1.ckt test2

.print op v(nodes) v2(r3)
.op
.list
.end
