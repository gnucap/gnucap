* nor-test
V2 1 0 10V
V1 4 0 10V
U2 2 0 4 4 3 5 CMOS NOR
V3 5 0 10V
U1 3 0 4 4 1 2 CMOS NOR
.model CMOS LOGIC
.print dc V(V2) V(V3) V(U1) V(U2) logic(u*)
.dc V2 0 10 2
.status notime
.END
