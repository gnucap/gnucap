This is the title
*this is a comment
VIN 12 0 AC .5
EIN 0 9 12 0 1
M1 3 9 10 11 MOD1 W=59U L=10U
M2 4 12 10 11 MOD1 W=59U L=10U
M3 3 3 1 1 MOD2 W=8U L=10U
M4 4 3 1 1 MOD2 W=8U L=10U
M5 10 8 11 11 MOD1 W=51U L=10U
M6 5 4 1 1 MOD2 W=39U L=10U
M7 5 8 11 11 MOD1 W=949U L=10U
M8 8 8 11 11 MOD1 W=56U L=10U
IREF 1 8 10U
*M9 8 8 7 1 MOD2 W=10U L=10U
*M10 7 7 6 1 MOD2 W=11U L=10U
*M11 6 6 1 1 MOD2 W=10U L=10U
.MODEL MOD1 NMOS Level=2 VTO=1.0 KP=17U GAMMA=1.3 LAMBDA=0.01 PHI=0.7
.MODEL MOD2 PMOS Level=2 VTO=-1.0 KP=8U GAMMA=0.6 LAMBDA=0.02 PHI=0.6
CC 4 5 6PF
VCC 1 0 DC +5
VSS 11 0 DC -5
*.AC DEC 10 1HZ 20M
*.plot ac vdb(5) vp(5)
*>.options out=200 vmin=-5.5 vmax=5.5 dampstrategy=2
*>.print op v(1 3 4 5 8 9 10 11 12)
.op trace iterations
*>.stat notime
.END
