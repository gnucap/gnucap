# HSPICE style PWL, out of order, bogus answers
v1 1 0 dc 1 ac 1
r1 1 2 1k
r2 2 0 1k
e1 3 0 2 0 PWL(1) 0,0 1,1 4,2 9,3 160,4 25,5
r3 3 0 10k
.list
.print op v(1) v(2) v(3)
.op
.print dc v(nodes)
.dc v1 -10 10 1
.dc v1 1 1000 decade 5
.dc v1 32 68 9
.end
