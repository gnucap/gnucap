difpair ckt - simple differential pair
* modified from Spice-3 examples

*>.opt rstray cstray
*.tf v(5) vin
*.dc vin -0.25 0.25 0.005

vin 1 0 sin(0 0.1 5meg) ac 1 dc 0
vcc 8 0 12
vee 9 0 -12
q1 4 2 6 0 qnl
q2 5 3 6 0 qnl
rs1 1 2 1k
rs2 3 0 1k
rc1 4 8 10k
rc2 5 8 10k
q3 6 7 9 0 qnl
q4 7 7 9 0 qnl
rbias 7 8 20k
*.model qnl npn(bf=80 rb=100 ccs=2pf tf=0.3ns tr=6ns cje=3pf cjc=2pf
*+   va=50)
.model qnl npn(bf=80 rb=100 va=50 ccs=20pf)

*>.print tran v(4) v(5)
*>.print op ccs(q*)
.op
.plot tran v(5)
*>.plot tran v(5)(4,8)
.tran 5ns 500ns
*>.print tran qcs(q*)
*>.tran 5ns 500ns
*>.print tran ccs(q*)
*>.tran 5ns 500ns
*>.print tran vcs(q*)
*>.tran 5ns 500ns

.plot ac vm(5) vp(5)
*>.plot ac vm(5)(-70,90) vp(5)(-70,90)
.ac dec 10 1 10ghz

.end
