A 1153 node circuit
Vin 1 0 dc 1 ac 1
x1 1 2 0 eq32
.subckt eq32 1 3 g
x1 1 2 g eq16
x2 2 3 g eq16
.ends eq32
.subckt eq16 1 5 g
x1 1 2 g eq4
x2 2 3 g eq4
x3 3 4 g eq4
x4 4 5 g eq4
.ends eq16
.subckt eq4 1 5 g
x1 1 2 g eq
x2 2 3 g eq
x3 3 4 g eq
x4 4 5 g eq
.ends eq4
.subckt eq 31 37 g
R101a   35   1  50.K
R101b   36   1  50.K
R102a   32   4  50.K
R102b   33   4  50.K
R103a   35   7  50.K
R103b   36   7  50.K
R104a   32  10  50.K
R104b   33  10  50.K
R105a   35  13  50.K
R105b   36  13  50.K
R106a   32  16  50.K
R106b   33  16  50.K
R107a   35  19  50.K
R107b   36  19  50.K
R108a   32  22  50.K
R108b   33  22  50.K
R109a   35  25  50.K
R109b   36  25  50.K
R110a   32  28  50.K
R110b   33  28  50.K
C1      1   2  1.5u
C2      4   5  748.n
C3      7   8  408.n
C4     10  11  206.n
C5     13  14  100.n
C6     16  17  50.9n
C7     19  20  25.3n
C8     22  23  12.7n
C9     25  26  5.9n
C10    28  29  2.95n
C11     2   3  15.n
C12     5   6  6.8n
C13     8   9  3.3n
C14    11  12  1.8n
C15    14  15  1.n
C16    17  18  470.p
C17    20  21  220.p
C18    23  24  120.p
C19    26  27  68.p
C20    29  30  33.p
R1      3   g  475.K
R2      6   g  536.K
R3      9   g  549.K
R4     12   g  499.K
R5     15   g  464.K
R6     18   g  475.K
R7     21   g  523.K
R8     24   g  475.K
R9     27   g  412.K
R10    30   g  422.K
G5a     2   g   3   g   -.000416666
R11     2   g  2.4K
G5b     5   g   6   g   -.000416666
R12     5   g  2.4K
G6a     8   g   9   g   -.000454545
R13     8   g  2.2K
G6b    11   g  12   g   -.000454545
R14    11   g  2.2K
G7a    14   g  15   g   -.000454545
R15    14   g  2.2K
G7b    17   g  18   g   -.000454545
R16    17   g  2.2K
G8a    20   g  21   g   -.000454545
R17    20   g  2.2K
G8b    23   g  24   g   -.000454545
R18    23   g  2.2K
G9a    26   g  27   g   -.000416666
R19    26   g  2.4K
G9b    29   g  30   g   -.000416666
R20    29   g  2.4K
R29    31  32  9.1K
R30    33  34  9.1K
R31    34  35  9.1K
R32    36  37  9.1K
C25    31  32  150.p
C26    33  34  150.p
C27    34  35  150.p
C28    36  37  150.p
E2     34   g  32  33  10.K
E3     37   g  35  36  10.K
.ends eq
.print op iter(0) v(1) v(2)
.print dc v(2)
.print ac vm(2) vdb(2) vp(2)
.dc Vin 1 10 1
.ac oct 1 31.25 16000
.end
