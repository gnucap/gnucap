' exp test, periodic
.option out=170 list
.param ppp=50n
.subckt esource (a b)
*.parameter p
v1 (a b) exp  iv= 0.  pv= 1.  td1=p/20  tau1=p/4  td2=p/2  tau2=p/4  period=p
.ends
x1 (1 0) esource p=ppp
*x2 (2 0) esource p=20n
.print tran v(1)
.param ppp=20n
.tran 0 100n 100n trace all
.param ppp=50n
.tran  trace all
.list
*>.status notime
.end
