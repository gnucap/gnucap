'
V1  1  0  DC   1.
E1  2  0  1  0  TANH  gain= 100.  limit= 0.01
.print dc v nodes
.dc v1 -.00000001 .00000001 .000000001
.dc v1 -.0000001 .0000001 .00000001
.dc v1 -.000001 .000001 .0000001
.dc v1 -.00001 .00001 .000001
.dc v1 -.0001 .0001 .00001
.dc v1 -.001 .001 .0001
.dc v1 -.01 .01 .001
.dc v1 -.1 .1 .01
.dc v1 -1 1 .1
.dc v1 -10 10 1
.dc v1 -100 100 10
.dc v1 -1000 1000 100
.dc v1 -10k 10k 1k
.dc v1 -100k 100k 10k
.dc v1 -1000k 1000k 100k
.dc v1 -10000k 10000k 1000k
.end
