' a test of the delete command
V1 1 0 1
R1 1 2 1
R2 2 0 1
R31 2 3 1
R32 3 0 2
L 3 4 5
C1 4 0 5
C2 4 5 5
C3 5 0 2
.option trace
.print op v(nodes)
.list
.op
.delete L
.list
.op
.delete R3*
.list
.op
.delete L*
.list
.op
.delete c*
.list
.op
.delete r2
.list
.op
.delete r*
.list
.op
.end
