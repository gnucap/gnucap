'
V1   1  0  dc 1. ac 9
X1   1  2  3  4  5  6  7  8  9  zzzz
.subckt zzzz  9  8  7  6  5  4  3  2  1 
R1   1  0  1.
R2   1  2  1.
R3   2  3  1.
R4   3  4  1.
R5   4  5  1.
R6   5  6  1.
R7   6  7  1.
R8   7  8  1.
R9   8  9  1.
R10   9  0  1.
.ends
.print op v nodes
.op
.print ac v nodes
.ac 1k
*>.status notime
.end
