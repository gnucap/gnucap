#Transmission lines

.width out=160

V1 1 0 gen(1)

# matched
R1s 1 11 50
T1 11 0 12 0 z=50 f=10meg nl=.25
R1l 12 0 50

# open stub
R2s 1 21 50
T2 21 0 22 0 z=50 f=10meg nl=.25
R2l 22 0 1e99

# shorted stub
R3s 1 31 50
T3 31 0 32 0 z=50 f=10meg nl=.25
R3l 32 0 .001

# lo-z load
R4s 1 41 50
T4 41 0 42 0 z=50 f=10meg nl=.25
R4l 42 0 25

# hi-z load
R5s 1 51 50
T5 51 0 52 0 z=50 f=10meg nl=.25
R5l 52 0 100

.list
.print ac v nodes

# nominal-z drive
.ac 0 40meg 2meg

# very lo-z drive
.modify R?s=.1
.ac

# slightly lo-z drive
.modify R?s=25
.ac

# hi-z drive
.modify R?s=100
.ac

.end

