
.param p1  = '1/(8.854e-12*3.9)'

v1 1 0 dc 'p1'
v2 2 0 dc '1/(8.854e-12*3.9)'
v3 3 0 dc '1/8.854e-12/3.9'  
v4 4 0 dc '8.854e-12*3.9'
v5 5 0 dc '8.854e-12'
v6 6 0 dc '1.e-12'
v7 7 0 dc  1.e-12

.print op v(1) v(2) v(3) v(4) v(5) v(6) v(7)
.op 

.end
