'c check
.option short=.1u
v1 1 0  pulse(0 1 0 .0001 .0001 1k 1k) ac 1
r1 1 2 .01
c2 2 0 1
.list
.print tran v(1) v(2)
.tran .001 .01 0
.tran .01 .10 0
.tran .1 1 0
.tran 1 10 0
.status notime
.end
