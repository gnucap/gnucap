
.get d_cccs.1.ckt
.print ac v(1)
.ac
.end
