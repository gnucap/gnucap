
u1 1 2 3 4 5 mos nand
.model mos nmos
.op
.end
