# semiconductor "resistor" test
.param pw=2u pl=1u
v1 1 0 dc 2 ac 5
r1 1 2 1k
r2 2 0 t1 (w=pw l=pl)
.model t1 r rsh=1k
.print op v(nodes) r(r*)
.print ac v(nodes) 
.op
.ac
.list
.end
