* switch as negative resistance oscillator
* Spice netlister for gnetlist
SW1 1 0 1 0 SWITCH1
C1 1 0 1n
I1 0 1 100u
.MODEL SWITCH1 SW VT=2.5 VH=2.475 RON=1 ROFF=10MEG
.print tran V(1)
*>.print tran + r(SW1) iter(0) input(sw1) timef(sw1) control(0)
.option method=trap itl6=0
.tran 10e-6 200e-6  trace iter
*>.status notime
.END
